* SPICE3 file created from XNOR2IN.ext - technology: scmos

.include TSMC_180nm.txt
.option scale=0.09u

.param SUPPLY = 1.8
.global gnd

Vdd vdd gnd 'SUPPLY'

V_in_a vin1 gnd PULSE(1.8 0 0ns 100ps 100ps 20ns 40ns)
V_in_b vin2 gnd PULSE(1.8 0 0ns 100ps 100ps 40ns 80ns)

M1000 XOR2IN_0/NAND2IN_0/a_n1_n23# vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=100 ps=90
M1001 XOR2IN_0/NAND2IN_2/vin2 vin1 vdd XOR2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=190 ps=166
M1002 XOR2IN_0/NAND2IN_2/vin2 vin2 XOR2IN_0/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1003 XOR2IN_0/NAND2IN_2/vin2 vin2 vdd XOR2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 XOR2IN_0/NAND2IN_1/a_n1_n23# vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1005 XOR2IN_0/NAND2IN_3/vin1 vin1 vdd XOR2IN_0/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1006 XOR2IN_0/NAND2IN_3/vin1 XOR2IN_0/NAND2IN_2/vin2 XOR2IN_0/NAND2IN_1/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1007 XOR2IN_0/NAND2IN_3/vin1 XOR2IN_0/NAND2IN_2/vin2 vdd XOR2IN_0/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 XOR2IN_0/NAND2IN_2/a_n1_n23# vin2 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1009 XOR2IN_0/NAND2IN_3/vin2 vin2 vdd XOR2IN_0/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1010 XOR2IN_0/NAND2IN_3/vin2 XOR2IN_0/NAND2IN_2/vin2 XOR2IN_0/NAND2IN_2/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1011 XOR2IN_0/NAND2IN_3/vin2 XOR2IN_0/NAND2IN_2/vin2 vdd XOR2IN_0/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1012 XOR2IN_0/NAND2IN_3/a_n1_n23# XOR2IN_0/NAND2IN_3/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1013 NOT_0/in XOR2IN_0/NAND2IN_3/vin1 vdd XOR2IN_0/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1014 NOT_0/in XOR2IN_0/NAND2IN_3/vin2 XOR2IN_0/NAND2IN_3/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1015 NOT_0/in XOR2IN_0/NAND2IN_3/vin2 vdd XOR2IN_0/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1016 vout NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1017 vout NOT_0/in vdd NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
C0 XOR2IN_0/NAND2IN_2/vin2 vin2 0.39fF
C1 NOT_0/in XOR2IN_0/NAND2IN_3/vin2 0.06fF
C2 XOR2IN_0/NAND2IN_3/w_n16_n4# XOR2IN_0/NAND2IN_3/vin2 0.10fF
C3 XOR2IN_0/NAND2IN_3/vin1 XOR2IN_0/NAND2IN_2/vin2 0.06fF
C4 vdd gnd 0.11fF
C5 XOR2IN_0/NAND2IN_2/vin2 gnd 0.19fF
C6 NOT_0/w_n7_n3# NOT_0/in 0.07fF
C7 vin1 XOR2IN_0/NAND2IN_1/w_n16_n4# 0.10fF
C8 vout gnd 0.07fF
C9 gnd vin2 0.09fF
C10 XOR2IN_0/NAND2IN_2/w_n16_n4# vdd 0.11fF
C11 XOR2IN_0/NAND2IN_3/vin1 gnd 0.13fF
C12 vdd vin1 0.06fF
C13 XOR2IN_0/NAND2IN_2/w_n16_n4# XOR2IN_0/NAND2IN_2/vin2 0.10fF
C14 vdd XOR2IN_0/NAND2IN_0/w_n16_n4# 0.11fF
C15 vdd NOT_0/in 0.08fF
C16 vdd XOR2IN_0/NAND2IN_3/w_n16_n4# 0.11fF
C17 XOR2IN_0/NAND2IN_2/w_n16_n4# vin2 0.10fF
C18 XOR2IN_0/NAND2IN_2/vin2 XOR2IN_0/NAND2IN_0/w_n16_n4# 0.08fF
C19 vdd XOR2IN_0/NAND2IN_3/vin2 0.08fF
C20 vin2 XOR2IN_0/NAND2IN_0/w_n16_n4# 0.10fF
C21 XOR2IN_0/NAND2IN_3/vin2 XOR2IN_0/NAND2IN_2/vin2 0.06fF
C22 XOR2IN_0/NAND2IN_3/vin1 XOR2IN_0/NAND2IN_3/w_n16_n4# 0.10fF
C23 vin1 gnd 0.27fF
C24 vdd NOT_0/w_n7_n3# 0.06fF
C25 NOT_0/in gnd 0.01fF
C26 vdd XOR2IN_0/NAND2IN_1/w_n16_n4# 0.11fF
C27 vout NOT_0/w_n7_n3# 0.03fF
C28 XOR2IN_0/NAND2IN_3/vin2 gnd 0.06fF
C29 XOR2IN_0/NAND2IN_2/vin2 XOR2IN_0/NAND2IN_1/w_n16_n4# 0.10fF
C30 XOR2IN_0/NAND2IN_3/vin1 XOR2IN_0/NAND2IN_1/w_n16_n4# 0.08fF
C31 vdd XOR2IN_0/NAND2IN_2/vin2 0.08fF
C32 vin1 XOR2IN_0/NAND2IN_0/w_n16_n4# 0.10fF
C33 vdd vout 0.06fF
C34 XOR2IN_0/NAND2IN_2/w_n16_n4# XOR2IN_0/NAND2IN_3/vin2 0.08fF
C35 NOT_0/in XOR2IN_0/NAND2IN_3/w_n16_n4# 0.08fF
C36 vdd XOR2IN_0/NAND2IN_3/vin1 0.43fF
C37 vout Gnd 0.09fF
C38 NOT_0/w_n7_n3# Gnd 0.61fF
C39 vdd Gnd 0.81fF
C40 NOT_0/in Gnd 0.38fF
C41 XOR2IN_0/NAND2IN_3/vin1 Gnd 0.54fF
C42 XOR2IN_0/NAND2IN_3/w_n16_n4# Gnd 1.16fF
C43 XOR2IN_0/NAND2IN_3/vin2 Gnd 0.55fF
C44 XOR2IN_0/NAND2IN_2/vin2 Gnd 0.80fF
C45 XOR2IN_0/NAND2IN_2/w_n16_n4# Gnd 1.16fF
C46 XOR2IN_0/NAND2IN_1/w_n16_n4# Gnd 1.16fF
C47 vin2 Gnd 1.17fF
C48 vin1 Gnd 2.31fF
C49 XOR2IN_0/NAND2IN_0/w_n16_n4# Gnd 1.16fF

.tran 1n 600n

.control
run
set color0 = rgb:f/f/e
set color1 = black
plot v(vin1) v(vin2)+2 (vout)+4
hardcopy image.ps v(vin1) v(vin2)+2 (vout)+4
.end
.endc