Testbench for all individual components

.include TSMC_180nm.txt
.include All_Gates.sub
.include And.sub
.include Enable.sub
.include Decoder.sub
.include AdderSubtractor.sub
.include Comparator.sub
.include ALU.sub


.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd node_x gnd 'SUPPLY'

V_in_a3 node_a3 gnd PULSE(0 1.8 0ns 100ps 100ps 10ns 50ns)
V_in_b3 node_b3 gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 70ns)
V_in_a2 node_a2 gnd PULSE(0 1.8 0ns 100ps 100ps 30ns 70ns)
V_in_b2 node_b2 gnd PULSE(0 1.8 0ns 100ps 100ps 40ns 50ns)
V_in_a1 node_a1 gnd PULSE(0 1.8 0ns 100ps 100ps 40ns 70ns)
V_in_b1 node_b1 gnd PULSE(0 1.8 0ns 100ps 100ps 30ns 50ns)
V_in_a0 node_a0 gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 50ns)
V_in_b0 node_b0 gnd PULSE(0 1.8 0ns 100ps 100ps 10ns 70ns)

* ----------------------------------And Test-----------------------------------------------

* X_AND node_out3 node_out2 node_out1 node_out0 node_a3 node_a2 node_a1 node_a0 node_b3 node_b2 node_b1 node_b0 node_x gnd And

* C1 node_out0 gnd 100f
* C2 node_out1 gnd 100f
* C3 node_out2 gnd 100f
* C4 node_out3 gnd 100f


* .tran 1n 800n

* .control
* run
* set color0 = rgb:f/f/e
* set color1 = black
* plot v(node_a0) v(node_b0)+2 v(node_out0)+4 v(node_a1)+6 v(node_b1)+8 v(node_out1)+10 v(node_a2)+12 v(node_b2)+14 v(node_out2)+16 v(node_a3)+18 v(node_b3)+20 v(node_out3)+22

* hardcopy image.ps v(node_a0) v(node_b0)+2 v(node_out0)+4 v(node_a1)+6 v(node_b1)+8 v(node_out1)+10 v(node_a2)+12 v(node_b2)+14 v(node_out2)+16 v(node_a3)+18 v(node_b3)+20 v(node_out3)+22
* .end
* .endc

* ------------------------------------comparator test--------------------------------------

* V_in_en node_en gnd PULSE(0 1.8 0ns 100ps 100ps 800ns 1000ns)

* X_Comp Greater Equal Less node_a3 node_a2 node_a1 node_a0 node_b3 node_b2 node_b1 node_b0 node_en node_x gnd Comparator

* C1 Greater gnd 100f
* C2 Equal gnd 100f
* C3 Less gnd 100f

* .tran 1n 800n

* .control
* run
* set color0 = rgb:f/f/e
* set color1 = black
* plot v(node_a0) v(node_b0)+8 v(node_a1)+2 v(node_b1)+10 v(node_a2)+4 v(node_b2)+12 v(node_a3)+6 v(node_b3)+14 v(Greater)+16 v(Equal)+18 v(Less)+20

* hardcopy image.ps v(node_a0) v(node_b0)+8 v(node_a1)+2 v(node_b1)+10 v(node_a2)+4 v(node_b2)+12 v(node_a3)+6 v(node_b3)+14 v(Greater)+16 v(Equal)+18 v(Less)+20

* .end
* .endc

* -----------------------------------Adder Subtractor Test---------------------------------
* V_in_en node_M gnd PULSE(1.8 0 0ns 100ps 100ps 400ns 800ns)

* X_add node_out3 node_out2 node_out1 node_out0 Carry node_a3 node_a2 node_a1 node_a0 node_b3 node_b2 node_b1 node_b0 node_M node_x gnd AdderSubtractor


* C1 node_out0 gnd 100f
* C2 node_out1 gnd 100f
* C3 node_out2 gnd 100f
* C4 node_out3 gnd 100f
* C5 Carry gnd 100f

* .tran 1n 800n

* .control
* run
* set color0 = rgb:f/f/e
* set color1 = black
* plot  v(node_M)-2 v(node_a0) v(node_b0)+2 v(node_out0)+4 v(node_a1)+6 v(node_b1)+8 v(node_out1)+10 v(node_a2)+12 v(node_b2)+14 v(node_out2)+16 v(node_a3)+18 v(node_b3)+20 v(node_out3)+22 v(Carry)+24

* hardcopy image.ps v(node_M)-2 v(node_a0) v(node_b0)+2 v(node_out0)+4 v(node_a1)+6 v(node_b1)+8 v(node_out1)+10 v(node_a2)+12 v(node_b2)+14 v(node_out2)+16 v(node_a3)+18 v(node_b3)+20 v(node_out3)+22
* .end
* .endc

* -----------------------------------ALU Test------------------------------------------
V_in_s1 Sel1 gnd PULSE(1.8 0 0ns 100ps 100ps 400ns 800ns)
V_in_s0 Sel0 gnd PULSE(1.8 0 0ns 100ps 100ps 200ns 400ns)

X_ALU CarryOut node_out3 node_out2 node_out1 node_out0 node_a3 node_a2 node_a1 node_a0 node_b3 node_b2 node_b1 node_b0 Sel1 Sel0 node_x gnd ALU


C1 node_out0 gnd 100f
C2 node_out1 gnd 100f
C3 node_out2 gnd 100f
C4 node_out3 gnd 100f
C5 CarryOut gnd 100f

.tran 1n 800n

.control
run
set color0 = rgb:f/f/e
set color1 = black
plot v(Sel0)-4 v(Sel1)-2 v(node_a0) v(node_b0)+2 v(node_out0)+4 v(node_a1)+6 v(node_b1)+8 v(node_out1)+10 v(node_a2)+12 v(node_b2)+14 v(node_out2)+16 v(node_a3)+18 v(node_b3)+20 v(node_out3)+22 v(CarryOut)+24

hardcopy image.ps v(Sel0)-4 v(Sel1)-2 v(node_a0) v(node_b0)+2 v(node_out0)+4 v(node_a1)+6 v(node_b1)+8 v(node_out1)+10 v(node_a2)+12 v(node_b2)+14 v(node_out2)+16 v(node_a3)+18 v(node_b3)+20 v(node_out3)+22 v(CarryOut)+24
.end
.endc

* ------------------------------------------Decoder Test---------------------------------------------
* V_in_s1 Sel1 gnd PULSE(1.8 0 0ns 100ps 100ps 400ns 800ns)
* V_in_s0 Sel0 gnd PULSE(1.8 0 0ns 100ps 100ps 200ns 400ns)

* X_Decoder node_out3 node_out2 node_out1 node_out0 Sel1 Sel0 node_x gnd Decoder


* C1 node_out0 gnd 100f
* C2 node_out1 gnd 100f
* C3 node_out2 gnd 100f
* C4 node_out3 gnd 100f

* .tran 1n 800n

* .control
* run
* set color0 = rgb:f/f/e
* set color1 = black
* plot v(Sel0) v(Sel1)+2 v(node_out0)+4 v(node_out1)+6 v(node_out2)+8 v(node_out3)+10
* hardcopy image.ps v(Sel0) v(Sel1)+2 v(node_out0)+4 v(node_out1)+6 v(node_out2)+8 v(node_out3)+10

* .end
* .endc

* --------------------------- Enable -----------------------------
* V_in_en node_M gnd PULSE(1.8 0 0ns 100ps 100ps 400ns 800ns)

* X_Enable node_aout3 node_aout2 node_aout1 node_aout0 node_out3 node_out2 node_out1 node_out0 node_a3 node_a2 node_a1 node_a0 node_b3 node_b2 node_b1 node_b0 node_M node_x gnd Enable

* C1 node_out0 gnd 100f
* C2 node_out1 gnd 100f
* C3 node_out2 gnd 100f
* C4 node_out3 gnd 100f

* .tran 1n 800n

* .control
* run
* set color0 = rgb:f/f/e
* set color1 = black
* plot  v(node_M)-2 v(node_a0) v(node_b0)+2 v(node_out0)+4 v(node_a1)+6 v(node_b1)+8 v(node_out1)+10 v(node_a2)+12 v(node_b2)+14 v(node_out2)+16 v(node_a3)+18 v(node_b3)+20 v(node_out3)+22 

* hardcopy image.ps v(node_M)-2 v(node_a0) v(node_b0)+2 v(node_out0)+4 v(node_a1)+6 v(node_b1)+8 v(node_out1)+10 v(node_a2)+12 v(node_b2)+14 v(node_out2)+16 v(node_a3)+18 v(node_b3)+20 v(node_out3)+22
* .end
* .endc