magic
tech scmos
timestamp 1699609590
<< metal1 >>
rect -843 -107 -744 -104
rect -596 -107 -416 -104
rect -748 -196 -745 -176
rect -526 -207 -511 -204
rect -198 -207 -178 -204
rect -884 -256 -861 -253
rect -856 -256 -838 -253
rect -748 -298 -745 -242
rect -514 -253 -511 -207
rect -527 -256 -511 -253
rect -884 -313 -838 -310
rect -841 -439 -838 -313
rect -814 -403 -811 -344
rect -748 -355 -745 -325
rect -699 -390 -646 -387
rect -814 -406 -788 -403
rect -776 -432 -773 -423
rect -782 -435 -773 -432
rect -757 -439 -754 -425
rect -841 -442 -754 -439
rect -886 -474 -859 -471
rect -740 -493 -737 -403
rect -649 -451 -646 -390
rect -527 -432 -524 -256
rect -514 -418 -511 -310
rect -420 -356 -328 -353
rect -241 -401 -178 -398
rect -401 -420 -398 -404
rect -401 -423 -338 -420
rect -486 -426 -463 -423
rect -447 -432 -444 -423
rect -527 -435 -444 -432
rect -337 -437 -333 -435
rect -313 -451 -309 -433
rect -649 -454 -309 -451
rect -780 -496 -700 -493
<< m2contact >>
rect -749 -201 -744 -196
rect -814 -231 -809 -226
rect -748 -242 -743 -237
rect -861 -257 -856 -252
rect -486 -231 -481 -226
rect -749 -303 -744 -298
rect -748 -325 -743 -320
rect -814 -344 -809 -339
rect -704 -365 -699 -360
rect -787 -435 -782 -430
rect -859 -475 -853 -469
rect -712 -407 -707 -402
rect -481 -357 -476 -352
rect -390 -391 -385 -386
rect -482 -407 -477 -402
rect -514 -423 -509 -418
rect -491 -426 -486 -421
rect -338 -442 -333 -437
<< metal2 >>
rect -860 -432 -857 -257
rect -814 -339 -811 -231
rect -748 -237 -745 -201
rect -748 -320 -745 -303
rect -486 -341 -483 -231
rect -809 -344 -483 -341
rect -489 -356 -481 -353
rect -489 -361 -486 -356
rect -699 -364 -486 -361
rect -707 -406 -482 -403
rect -514 -426 -491 -423
rect -860 -435 -787 -432
rect -514 -471 -511 -426
rect -388 -439 -385 -391
rect -388 -442 -338 -439
rect -853 -474 -511 -471
use XOR2IN  XOR2IN_1
timestamp 1698769192
transform 1 0 -408 0 1 -205
box -106 -118 213 101
use XOR2IN  XOR2IN_0
timestamp 1698769192
transform 1 0 -736 0 1 -205
box -106 -118 213 101
use AND2IN  AND2IN_0
timestamp 1698685374
transform 1 0 -789 0 1 -411
box -2 -15 94 58
use AND2IN  AND2IN_1
timestamp 1698685374
transform 1 0 -479 0 1 -411
box -2 -15 94 58
use OR2IN  OR2IN_0
timestamp 1698686464
transform 1 0 -316 0 1 -381
box -25 -54 77 28
<< labels >>
rlabel metal1 -828 -106 -827 -105 5 vdd
rlabel metal1 -883 -255 -882 -254 3 vin1
rlabel metal1 -882 -312 -881 -311 3 vin2
rlabel metal1 -184 -206 -183 -205 7 vout
rlabel metal1 -186 -400 -185 -399 1 vcout
rlabel metal1 -739 -495 -738 -494 1 gnd
rlabel metal1 -882 -473 -879 -472 1 vcin
<< end >>
