magic
tech scmos
timestamp 1699715518
<< metal1 >>
rect 647 1872 650 1926
rect 859 1874 862 1926
rect 1071 1876 1074 1926
rect 1134 1867 1179 1868
rect 924 1865 975 1867
rect 746 1863 762 1865
rect 518 1860 559 1863
rect 606 1862 762 1863
rect 821 1864 975 1865
rect 1029 1865 1179 1867
rect 1029 1864 1144 1865
rect 821 1862 929 1864
rect 606 1860 749 1862
rect 294 1753 500 1756
rect 294 1727 297 1753
rect 518 1692 521 1860
rect 647 1815 650 1850
rect 859 1817 862 1852
rect 1071 1819 1074 1854
rect 1262 1820 1265 1926
rect 1293 1876 2654 1879
rect 621 1799 756 1802
rect 839 1801 967 1804
rect 1054 1803 1166 1806
rect 538 1793 544 1796
rect 545 1756 549 1785
rect 538 1753 549 1756
rect 561 1751 565 1782
rect 579 1774 583 1783
rect 561 1748 735 1751
rect 757 1732 761 1785
rect 773 1758 777 1786
rect 791 1783 908 1786
rect 969 1738 973 1787
rect 985 1767 989 1787
rect 1003 1785 1107 1788
rect 1293 1789 1296 1876
rect 2651 1859 2654 1876
rect 1167 1745 1171 1787
rect 1191 1786 1296 1789
rect 1167 1742 2684 1745
rect 969 1735 1884 1738
rect 757 1729 1088 1732
rect 1881 1728 1884 1735
rect 2681 1729 2684 1742
rect 2735 1729 2738 1926
rect 5099 1882 5638 1885
rect 2803 1876 5752 1879
rect 2803 1859 2806 1876
rect 2828 1748 4086 1751
rect 4083 1675 4086 1748
rect 4433 1685 4436 1753
rect 4640 1678 4643 1761
rect 2756 1519 3289 1522
rect 2602 1384 2838 1387
rect -953 1305 -505 1308
rect -953 262 -950 1305
rect 2835 1043 2838 1384
rect 5153 1135 5156 1272
rect 5409 1199 5412 1769
rect 5522 1199 5525 1748
rect 5638 1199 5641 1748
rect 5749 1198 5752 1876
rect 5153 1132 5305 1135
rect 2835 1040 3080 1043
rect -889 1020 -469 1023
rect -889 326 -886 1020
rect -435 590 -432 941
rect -418 610 -415 962
rect -398 627 -395 937
rect -380 643 -377 937
rect 9 650 12 938
rect 41 657 44 937
rect 67 664 70 935
rect 89 671 92 938
rect 2355 922 2358 941
rect 2940 907 2944 913
rect 553 904 2944 907
rect 89 668 526 671
rect 67 661 415 664
rect 41 654 299 657
rect 9 647 186 650
rect -380 640 45 643
rect -398 624 -66 627
rect -418 607 -182 610
rect -435 587 -295 590
rect -298 458 -295 587
rect -185 457 -182 607
rect -69 458 -66 624
rect 42 456 45 640
rect 183 456 186 647
rect 296 456 299 654
rect 412 458 415 661
rect 523 453 526 668
rect -546 434 -409 437
rect -546 310 -543 434
rect 553 420 556 904
rect 2990 900 2993 912
rect 691 897 2993 900
rect 691 456 694 897
rect 3011 892 3014 914
rect 804 889 3014 892
rect 804 458 807 889
rect 3034 884 3037 914
rect 920 881 3037 884
rect 920 455 923 881
rect 3056 876 3059 913
rect 1031 873 3059 876
rect 1031 456 1034 873
rect 3256 869 3259 912
rect 1172 866 3259 869
rect 1172 457 1175 866
rect 3274 861 3277 916
rect 1285 858 3277 861
rect 1285 455 1288 858
rect 3293 852 3296 912
rect 1401 849 3296 852
rect 1401 456 1404 849
rect 3313 844 3316 916
rect 1512 841 3316 844
rect 1512 458 1515 841
rect 5323 830 5326 1109
rect 5342 838 5345 1109
rect 1672 827 5326 830
rect 1672 456 1675 827
rect 5432 819 5435 1110
rect 5451 839 5454 1110
rect 1785 816 5435 819
rect 1785 456 1788 816
rect 5550 806 5553 1110
rect 5569 837 5572 1108
rect 1901 803 5553 806
rect 1901 456 1904 803
rect 5664 793 5667 1110
rect 2012 790 5667 793
rect 2012 457 2015 790
rect 2153 775 5340 778
rect 2153 456 2156 775
rect 2266 761 5449 764
rect 2266 458 2269 761
rect 2382 746 5567 749
rect 2382 457 2385 746
rect 5683 732 5686 1111
rect 2493 729 5686 732
rect 2493 456 2496 729
rect -828 307 -543 310
rect -820 281 -617 284
rect -1130 259 -918 262
rect -1130 162 -1127 259
rect -929 244 -911 247
rect -929 227 -926 244
rect -891 239 -887 248
rect -891 236 -774 239
rect -816 228 -813 236
rect -700 225 -697 253
rect -589 227 -586 238
rect -546 200 -543 307
rect -483 384 -412 387
rect 503 384 579 387
rect 1493 384 1569 387
rect -483 163 -480 384
rect -451 345 -415 348
rect -451 286 -448 345
rect -384 168 -381 348
rect -275 176 -272 348
rect -157 185 -154 348
rect -43 195 -40 348
rect 97 205 100 348
rect 206 215 209 348
rect 324 224 327 348
rect 438 233 441 348
rect 544 345 552 348
rect 557 345 574 348
rect -1130 159 -1080 162
rect -384 115 -381 163
rect -275 115 -272 171
rect -157 115 -154 180
rect -43 115 -40 190
rect 97 115 100 200
rect 206 115 209 210
rect 324 115 327 219
rect 438 115 441 228
rect 605 168 608 337
rect 714 176 717 346
rect 832 185 835 348
rect 946 195 949 348
rect 1086 205 1089 348
rect 1195 215 1198 348
rect 1313 224 1316 348
rect 1427 233 1430 348
rect 605 140 608 163
rect 714 150 717 171
rect 832 160 835 180
rect 946 171 949 190
rect 1086 182 1089 200
rect 1195 192 1198 210
rect 1313 204 1316 219
rect 1427 218 1430 228
rect 1586 140 1589 337
rect 1695 150 1698 337
rect 1813 160 1816 337
rect 1927 171 1930 337
rect 2067 182 2070 337
rect 2176 192 2179 337
rect 2294 204 2297 337
rect 2408 218 2411 337
rect -633 48 -630 65
rect -594 48 -591 65
<< m2contact >>
rect 646 1867 651 1872
rect 858 1869 863 1874
rect 1070 1871 1075 1876
rect 500 1752 505 1757
rect 646 1850 651 1855
rect 858 1852 863 1857
rect 1070 1854 1075 1859
rect 533 1792 538 1797
rect 533 1752 538 1757
rect 578 1769 583 1774
rect 735 1746 740 1751
rect 908 1783 914 1788
rect 771 1752 777 1758
rect 1107 1785 1112 1790
rect 2650 1854 2655 1859
rect 5094 1882 5099 1887
rect 5638 1882 5643 1887
rect 2802 1854 2807 1859
rect 5407 1769 5412 1774
rect 4638 1761 4643 1766
rect 4431 1753 4436 1758
rect 2823 1746 2828 1751
rect 2754 1514 2759 1519
rect 2610 1426 2615 1431
rect -505 1304 -500 1309
rect -380 1304 -375 1309
rect 5097 1335 5102 1340
rect 5520 1748 5526 1754
rect 5637 1748 5642 1753
rect 5296 1182 5301 1187
rect 2353 917 2358 922
rect 482 433 487 438
rect 5341 833 5346 838
rect 5450 834 5455 839
rect 5568 832 5573 837
rect 5340 775 5345 780
rect 5449 761 5454 766
rect 5567 746 5572 751
rect 573 433 578 438
rect 1471 433 1476 438
rect 1554 433 1559 438
rect 552 415 557 420
rect -617 280 -612 285
rect -700 253 -695 258
rect -774 236 -769 241
rect -589 238 -584 243
rect -453 281 -448 286
rect 539 343 544 348
rect 552 344 557 349
rect 437 228 442 233
rect 323 219 328 224
rect 205 210 210 215
rect 96 200 101 205
rect -44 190 -39 195
rect -158 180 -153 185
rect -276 171 -271 176
rect -385 163 -380 168
rect -556 157 -551 162
rect -485 158 -480 163
rect 1553 344 1558 349
rect 1426 228 1431 233
rect 1312 219 1317 224
rect 1194 210 1199 215
rect 1085 200 1090 205
rect 945 190 950 195
rect 831 180 836 185
rect 713 171 718 176
rect 604 163 609 168
rect 1426 213 1431 218
rect 1312 199 1317 204
rect 1194 187 1199 192
rect 1085 177 1090 182
rect 945 166 950 171
rect 831 155 836 160
rect 713 145 718 150
rect 2407 213 2412 218
rect 2293 199 2298 204
rect 2175 187 2180 192
rect 2066 177 2071 182
rect 1926 166 1931 171
rect 1812 155 1817 160
rect 1694 145 1699 150
rect 604 135 609 140
rect 1585 135 1590 140
<< pdm12contact >>
rect 984 1762 989 1767
<< metal2 >>
rect 910 1902 5525 1905
rect 647 1855 650 1867
rect 859 1857 862 1869
rect -500 1793 533 1796
rect -500 1308 -497 1793
rect 910 1788 914 1902
rect 1109 1882 5094 1885
rect 1071 1859 1074 1871
rect 1109 1790 1112 1882
rect 2655 1855 2802 1858
rect 583 1771 5407 1774
rect 989 1763 4638 1766
rect 505 1753 533 1756
rect 777 1755 4431 1758
rect 777 1754 782 1755
rect 5522 1754 5525 1902
rect 737 1740 740 1746
rect 960 1748 2823 1751
rect 960 1740 963 1748
rect 5638 1753 5641 1882
rect 737 1737 963 1740
rect 2612 1514 2754 1517
rect 2612 1431 2615 1514
rect 5102 1336 5299 1339
rect -500 1305 -380 1308
rect 5296 1187 5299 1336
rect -772 917 2353 920
rect -772 241 -769 917
rect 5342 780 5345 833
rect 5451 766 5454 834
rect 5569 751 5572 832
rect 487 434 573 437
rect 1476 434 1554 437
rect 553 349 556 415
rect 1517 345 1553 348
rect -612 281 -453 284
rect 539 258 542 343
rect -695 255 542 258
rect 1517 243 1520 345
rect -584 240 1520 243
rect 442 229 1426 232
rect 328 220 1312 223
rect 210 211 1194 214
rect 1431 214 2407 217
rect 101 201 1085 204
rect 1317 200 2293 203
rect -39 191 945 194
rect 1199 188 2175 191
rect -153 181 831 184
rect 1090 178 2066 181
rect -271 172 713 175
rect -380 164 604 167
rect 950 167 1926 170
rect -551 158 -485 161
rect 836 156 1812 159
rect 718 146 1694 149
rect 609 136 1585 139
use OR2IN  OR2IN_0
timestamp 1698686464
transform 1 0 -894 0 1 301
box -25 -54 77 28
use Decoder  Decoder_0
timestamp 1699639768
transform 1 0 -1042 0 1 129
box -53 -67 506 101
use Enable  Enable_0
timestamp 1699634857
transform 1 0 -411 0 1 358
box -5 -23 937 103
use Enable  Enable_1
timestamp 1699634857
transform 1 0 578 0 1 358
box -5 -23 937 103
use Enable  Enable_2
timestamp 1699634857
transform 1 0 1559 0 1 358
box -5 -23 937 103
use AdderSubtractor  AdderSubtractor_0
timestamp 1699694653
transform 1 0 -411 0 1 1305
box -67 -370 3149 427
use Comparator  Comparator_0
timestamp 1699693233
transform 1 0 3015 0 1 1166
box -76 -256 2141 522
use AND4Bit  AND4Bit_0
timestamp 1699631834
transform 1 0 5308 0 1 1112
box -12 -6 444 89
use OR3IN  OR3IN_0
timestamp 1698685914
transform 1 0 566 0 1 1835
box -25 -54 84 28
use OR3IN  OR3IN_1
timestamp 1698685914
transform 1 0 778 0 1 1837
box -25 -54 84 28
use OR2IN  OR2IN_1
timestamp 1698686464
transform 1 0 1188 0 1 1840
box -25 -54 77 28
use OR3IN  OR3IN_2
timestamp 1698685914
transform 1 0 990 0 1 1839
box -25 -54 84 28
<< labels >>
rlabel metal1 -632 49 -631 50 1 vinSel1
rlabel metal1 -593 50 -592 51 1 vinSel0
rlabel metal1 -383 120 -382 121 1 vina0
rlabel metal1 -274 118 -273 119 1 vina1
rlabel metal1 -156 118 -155 119 1 vina2
rlabel metal1 -42 116 -41 117 1 vina3
rlabel metal1 98 117 99 118 1 vinb0
rlabel metal1 207 117 208 118 1 vinb1
rlabel metal1 325 118 326 119 1 vinb2
rlabel metal1 439 117 440 118 1 vinb3
rlabel metal1 648 1922 649 1923 5 vout0
rlabel metal1 860 1920 861 1921 1 vout1
rlabel metal1 1072 1922 1073 1923 5 vout2
rlabel metal1 1263 1923 1264 1924 5 vout3
rlabel metal1 2736 1922 2737 1923 5 vcout
rlabel metal1 -565 1306 -564 1307 1 gnd
rlabel metal1 -797 1021 -795 1022 1 vdd
<< end >>
