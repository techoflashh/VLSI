* SPICE3 file created from XNOR2IN.ext - technology: scmos

.include TSMC_180nm.txt
.option scale=0.09u

.param SUPPLY = 1.8
.global gnd

Vdd vdd gnd 'SUPPLY'

V_in_a vin1 gnd PULSE(1.8 0 0ns 100ps 100ps 20ns 40ns)
V_in_b vin2 gnd PULSE(1.8 0 0ns 100ps 100ps 40ns 80ns)


M1000 XOR2IN_0/NAND2IN_0/a_n1_n23# vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=100 ps=90
M1001 XOR2IN_0/NAND2IN_2/vin1 vin1 vdd XOR2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=190 ps=166
M1002 XOR2IN_0/NAND2IN_2/vin1 vin2 XOR2IN_0/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1003 XOR2IN_0/NAND2IN_2/vin1 vin2 vdd XOR2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 XOR2IN_0/NAND2IN_1/a_n1_n23# vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1005 XOR2IN_0/NAND2IN_3/vin1 vin1 vdd XOR2IN_0/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1006 XOR2IN_0/NAND2IN_3/vin1 XOR2IN_0/NAND2IN_2/vin1 XOR2IN_0/NAND2IN_1/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1007 XOR2IN_0/NAND2IN_3/vin1 XOR2IN_0/NAND2IN_2/vin1 vdd XOR2IN_0/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 XOR2IN_0/NAND2IN_2/a_n1_n23# XOR2IN_0/NAND2IN_2/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1009 XOR2IN_0/NAND2IN_3/vin2 XOR2IN_0/NAND2IN_2/vin1 vdd XOR2IN_0/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1010 XOR2IN_0/NAND2IN_3/vin2 vin2 XOR2IN_0/NAND2IN_2/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1011 XOR2IN_0/NAND2IN_3/vin2 vin2 vdd XOR2IN_0/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1012 XOR2IN_0/NAND2IN_3/a_n1_n23# XOR2IN_0/NAND2IN_3/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1013 NOT_0/in XOR2IN_0/NAND2IN_3/vin1 vdd XOR2IN_0/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1014 NOT_0/in XOR2IN_0/NAND2IN_3/vin2 XOR2IN_0/NAND2IN_3/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1015 NOT_0/in XOR2IN_0/NAND2IN_3/vin2 vdd XOR2IN_0/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1016 vout NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1017 vout NOT_0/in vdd NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0

C0 XOR2IN_0/NAND2IN_2/vin1 vdd 0.08fF
C1 XOR2IN_0/NAND2IN_3/vin2 XOR2IN_0/NAND2IN_3/w_n16_n4# 0.10fF
C2 XOR2IN_0/NAND2IN_3/vin2 NOT_0/in 0.06fF
C3 NOT_0/w_n7_n3# vout 0.03fF
C4 vdd vout 0.06fF
C5 NOT_0/in XOR2IN_0/NAND2IN_3/w_n16_n4# 0.08fF
C6 XOR2IN_0/NAND2IN_2/vin1 XOR2IN_0/NAND2IN_3/vin1 0.06fF
C7 XOR2IN_0/NAND2IN_1/w_n16_n4# XOR2IN_0/NAND2IN_2/vin1 0.10fF
C8 XOR2IN_0/NAND2IN_3/vin2 vdd 0.08fF
C9 vin2 XOR2IN_0/NAND2IN_2/w_n16_n4# 0.10fF
C10 vdd XOR2IN_0/NAND2IN_3/w_n16_n4# 0.11fF
C11 XOR2IN_0/NAND2IN_2/vin1 XOR2IN_0/NAND2IN_2/w_n16_n4# 0.10fF
C12 NOT_0/w_n7_n3# NOT_0/in 0.07fF
C13 vdd NOT_0/in 0.08fF
C14 XOR2IN_0/NAND2IN_2/vin1 vin2 0.41fF
C15 XOR2IN_0/NAND2IN_3/vin1 XOR2IN_0/NAND2IN_3/w_n16_n4# 0.10fF
C16 vout gnd 0.07fF
C17 vdd XOR2IN_0/NAND2IN_0/w_n16_n4# 0.11fF
C18 NOT_0/w_n7_n3# vdd 0.06fF
C19 XOR2IN_0/NAND2IN_3/vin2 XOR2IN_0/NAND2IN_2/w_n16_n4# 0.08fF
C20 vin1 XOR2IN_0/NAND2IN_0/w_n16_n4# 0.10fF
C21 XOR2IN_0/NAND2IN_3/vin2 vin2 0.06fF
C22 vdd XOR2IN_0/NAND2IN_3/vin1 0.08fF
C23 NOT_0/in gnd 0.01fF
C24 XOR2IN_0/NAND2IN_1/w_n16_n4# vdd 0.11fF
C25 XOR2IN_0/NAND2IN_1/w_n16_n4# XOR2IN_0/NAND2IN_3/vin1 0.08fF
C26 vdd XOR2IN_0/NAND2IN_2/w_n16_n4# 0.11fF
C27 vin2 XOR2IN_0/NAND2IN_0/w_n16_n4# 0.10fF
C28 vin1 XOR2IN_0/NAND2IN_1/w_n16_n4# 0.10fF
C29 XOR2IN_0/NAND2IN_2/vin1 XOR2IN_0/NAND2IN_0/w_n16_n4# 0.08fF
C30 vout Gnd 0.02fF
C31 NOT_0/in Gnd 0.34fF
C32 NOT_0/w_n7_n3# Gnd 0.61fF
C33 XOR2IN_0/NAND2IN_3/vin1 Gnd 0.49fF
C34 XOR2IN_0/NAND2IN_3/w_n16_n4# Gnd 1.16fF
C35 XOR2IN_0/NAND2IN_3/vin2 Gnd 0.49fF
C36 vdd Gnd 0.26fF
C37 XOR2IN_0/NAND2IN_2/w_n16_n4# Gnd 1.16fF
C38 XOR2IN_0/NAND2IN_1/w_n16_n4# Gnd 1.16fF
C39 gnd Gnd 0.30fF
C40 vin2 Gnd 1.12fF
C41 vin1 Gnd 1.16fF
C42 XOR2IN_0/NAND2IN_0/w_n16_n4# Gnd 1.16fF

.tran 1n 600n

.control
run
set color0 = rgb:f/f/e
set color1 = black
plot v(vin1) v(vin2)+2 (vout)+4
hardcopy image.ps v(vin1) v(vin2)+2 (vout)+4
.end
.endc

