Question No 3 MajorityFunction

*temperature

.include TSMC_180nm.txt
.include All_Gates.sub

.subckt MUX Out A3 A2 A1 A0 S1 S0 vdd gnd
    X1 S1c S1 vdd gnd NOT
    X2 S0c S0 vdd gnd NOT
    X3 Out0 A0 S1c S0c vdd gnd AND3IN
    X4 Out1 A1 S1c S0 vdd gnd AND3IN
    X5 Out2 A2 S1 S0c vdd gnd AND3IN
    X6 Out3 A3 S1 S0 vdd gnd AND3IN
    X7 Out Out0 Out1 Out2 Out3 vdd gnd OR4IN
.ends MUX

.subckt MajorityFunction Out A2 A1 A0 vdd gnd
    X1 Out vdd A0 A0 gnd A2 A1 vdd gnd MUX
.ends MajorityFunction

.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd vdd gnd 'SUPPLY'

*inputPulses

Xm node_out node_a2 node_a1 node_a0 vdd gnd MajorityFunction 

C1 node_out gnd 0.5f

.tran 1n 640n

*delay

.control
run
quit
.end
.endc