* SPICE3 file created from ALU.ext - technology: scmos

.option scale=0.09u
.include TSMC_180nm.txt

.param SUPPLY = 1.8

.global gnd

Vdd vdd gnd 'SUPPLY'

V_in_a3 vina3 gnd DC 1.8
V_in_a2 vina2 gnd DC 0
V_in_a1 vina1 gnd DC 0
V_in_a0 vina0 gnd DC 0

V_in_b3 vinb3 gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)
V_in_b2 vinb2 gnd PULSE(0 1.8 0ns 100ps 100ps 60ns 120ns)
V_in_b1 vinb1 gnd PULSE(0 1.8 0ns 100ps 100ps 60ns 120ns)
V_in_b0 vinb0 gnd PULSE(0 1.8 0ns 100ps 100ps 60ns 120ns)

V_in_Sel1 vinSel1 gnd DC 1.8
V_in_Sel0 vinSel0 gnd DC 0


M1000 Decoder_0/AND4Bit_0/AND2IN_0/NAND2IN_0/a_n1_n23# Decoder_0/NOT_1/out gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=4083 ps=3675
M1001 Decoder_0/AND4Bit_0/AND2IN_0/NOT_0/in Decoder_0/NOT_1/out vdd Decoder_0/AND4Bit_0/AND2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=7215 ps=5837
M1002 Decoder_0/AND4Bit_0/AND2IN_0/NOT_0/in Decoder_0/NOT_0/out Decoder_0/AND4Bit_0/AND2IN_0/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1003 Decoder_0/AND4Bit_0/AND2IN_0/NOT_0/in Decoder_0/NOT_0/out vdd Decoder_0/AND4Bit_0/AND2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 OR2IN_0/vin1 Decoder_0/AND4Bit_0/AND2IN_0/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1005 OR2IN_0/vin1 Decoder_0/AND4Bit_0/AND2IN_0/NOT_0/in vdd Decoder_0/AND4Bit_0/AND2IN_0/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1006 Decoder_0/AND4Bit_0/AND2IN_1/NAND2IN_0/a_n1_n23# vinSel0 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1007 Decoder_0/AND4Bit_0/AND2IN_1/NOT_0/in vinSel0 vdd Decoder_0/AND4Bit_0/AND2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1008 Decoder_0/AND4Bit_0/AND2IN_1/NOT_0/in Decoder_0/NOT_0/out Decoder_0/AND4Bit_0/AND2IN_1/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1009 Decoder_0/AND4Bit_0/AND2IN_1/NOT_0/in Decoder_0/NOT_0/out vdd Decoder_0/AND4Bit_0/AND2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1010 OR2IN_0/vin2 Decoder_0/AND4Bit_0/AND2IN_1/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1011 OR2IN_0/vin2 Decoder_0/AND4Bit_0/AND2IN_1/NOT_0/in vdd Decoder_0/AND4Bit_0/AND2IN_1/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1012 Decoder_0/AND4Bit_0/AND2IN_2/NAND2IN_0/a_n1_n23# Decoder_0/NOT_1/out gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1013 Decoder_0/AND4Bit_0/AND2IN_2/NOT_0/in Decoder_0/NOT_1/out vdd Decoder_0/AND4Bit_0/AND2IN_2/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1014 Decoder_0/AND4Bit_0/AND2IN_2/NOT_0/in vinSel1 Decoder_0/AND4Bit_0/AND2IN_2/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1015 Decoder_0/AND4Bit_0/AND2IN_2/NOT_0/in vinSel1 vdd Decoder_0/AND4Bit_0/AND2IN_2/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1016 Enable_1/vinEn Decoder_0/AND4Bit_0/AND2IN_2/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1017 Enable_1/vinEn Decoder_0/AND4Bit_0/AND2IN_2/NOT_0/in vdd Decoder_0/AND4Bit_0/AND2IN_2/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1018 Decoder_0/AND4Bit_0/AND2IN_3/NAND2IN_0/a_n1_n23# vinSel0 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1019 Decoder_0/AND4Bit_0/AND2IN_3/NOT_0/in vinSel0 vdd Decoder_0/AND4Bit_0/AND2IN_3/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1020 Decoder_0/AND4Bit_0/AND2IN_3/NOT_0/in vinSel1 Decoder_0/AND4Bit_0/AND2IN_3/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1021 Decoder_0/AND4Bit_0/AND2IN_3/NOT_0/in vinSel1 vdd Decoder_0/AND4Bit_0/AND2IN_3/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1022 Enable_2/vinEn Decoder_0/AND4Bit_0/AND2IN_3/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1023 Enable_2/vinEn Decoder_0/AND4Bit_0/AND2IN_3/NOT_0/in vdd Decoder_0/AND4Bit_0/AND2IN_3/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1024 Decoder_0/NOT_1/out vinSel0 gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1025 Decoder_0/NOT_1/out vinSel0 vdd Decoder_0/NOT_1/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1026 Decoder_0/NOT_0/out vinSel1 gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1027 Decoder_0/NOT_0/out vinSel1 vdd Decoder_0/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1028 vout0 OR3IN_0/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1029 vout0 OR3IN_0/NOT_0/in vdd OR3IN_0/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1030 OR3IN_0/a_6_1# OR3IN_0/vin2 OR3IN_0/a_0_1# OR3IN_0/w_n19_n9# CMOSP w=12 l=2
+  ad=48 pd=32 as=48 ps=32
M1031 OR3IN_0/a_0_1# OR3IN_0/vin1 vdd OR3IN_0/w_n19_n9# CMOSP w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1032 OR3IN_0/NOT_0/in OR3IN_0/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=84 pd=66 as=0 ps=0
M1033 OR3IN_0/NOT_0/in OR3IN_0/vin3 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1034 OR3IN_0/NOT_0/in OR3IN_0/vin3 OR3IN_0/a_6_1# OR3IN_0/w_n19_n9# CMOSP w=12 l=2
+  ad=108 pd=42 as=0 ps=0
M1035 OR3IN_0/NOT_0/in OR3IN_0/vin2 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1036 vout1 OR3IN_1/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1037 vout1 OR3IN_1/NOT_0/in vdd OR3IN_1/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1038 OR3IN_1/a_6_1# OR3IN_1/vin2 OR3IN_1/a_0_1# OR3IN_1/w_n19_n9# CMOSP w=12 l=2
+  ad=48 pd=32 as=48 ps=32
M1039 OR3IN_1/a_0_1# OR3IN_1/vin1 vdd OR3IN_1/w_n19_n9# CMOSP w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1040 OR3IN_1/NOT_0/in OR3IN_1/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=84 pd=66 as=0 ps=0
M1041 OR3IN_1/NOT_0/in OR3IN_1/vin3 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1042 OR3IN_1/NOT_0/in OR3IN_1/vin3 OR3IN_1/a_6_1# OR3IN_1/w_n19_n9# CMOSP w=12 l=2
+  ad=108 pd=42 as=0 ps=0
M1043 OR3IN_1/NOT_0/in OR3IN_1/vin2 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1044 vout2 OR3IN_2/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1045 vout2 OR3IN_2/NOT_0/in vdd OR3IN_2/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1046 OR3IN_2/a_6_1# OR3IN_2/vin2 OR3IN_2/a_0_1# OR3IN_2/w_n19_n9# CMOSP w=12 l=2
+  ad=48 pd=32 as=48 ps=32
M1047 OR3IN_2/a_0_1# OR3IN_2/vin1 vdd OR3IN_2/w_n19_n9# CMOSP w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1048 OR3IN_2/NOT_0/in OR3IN_2/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=84 pd=66 as=0 ps=0
M1049 OR3IN_2/NOT_0/in OR3IN_2/vin3 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1050 OR3IN_2/NOT_0/in OR3IN_2/vin3 OR3IN_2/a_6_1# OR3IN_2/w_n19_n9# CMOSP w=12 l=2
+  ad=108 pd=42 as=0 ps=0
M1051 OR3IN_2/NOT_0/in OR3IN_2/vin2 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1052 OR2IN_0/vout OR2IN_0/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1053 OR2IN_0/vout OR2IN_0/NOT_0/in vdd OR2IN_0/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1054 OR2IN_0/NOT_0/in OR2IN_0/vin2 OR2IN_0/a_0_1# OR2IN_0/w_n19_n9# CMOSP w=12 l=2
+  ad=72 pd=36 as=48 ps=32
M1055 OR2IN_0/NOT_0/in OR2IN_0/vin2 gnd Gnd CMOSN w=4 l=2
+  ad=60 pd=46 as=0 ps=0
M1056 OR2IN_0/a_0_1# OR2IN_0/vin1 vdd OR2IN_0/w_n19_n9# CMOSP w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1057 OR2IN_0/NOT_0/in OR2IN_0/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1058 vout3 OR2IN_1/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1059 vout3 OR2IN_1/NOT_0/in vdd OR2IN_1/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1060 OR2IN_1/NOT_0/in OR2IN_1/vin2 OR2IN_1/a_0_1# OR2IN_1/w_n19_n9# CMOSP w=12 l=2
+  ad=72 pd=36 as=48 ps=32
M1061 OR2IN_1/NOT_0/in OR2IN_1/vin2 gnd Gnd CMOSN w=4 l=2
+  ad=60 pd=46 as=0 ps=0
M1062 OR2IN_1/a_0_1# OR2IN_1/vin1 vdd OR2IN_1/w_n19_n9# CMOSP w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1063 OR2IN_1/NOT_0/in OR2IN_1/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1064 Comparator_0/NOT_5/out Comparator_0/NOT_5/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1065 Comparator_0/NOT_5/out Comparator_0/NOT_5/in vdd Comparator_0/NOT_5/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1066 Comparator_0/NOT_6/out Comparator_0/NOT_6/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1067 Comparator_0/NOT_6/out Comparator_0/NOT_6/in vdd Comparator_0/NOT_6/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1068 Comparator_0/NOT_7/out Comparator_0/NOT_7/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1069 Comparator_0/NOT_7/out Comparator_0/NOT_7/in vdd Comparator_0/NOT_7/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1070 Comparator_0/OR4IN_0/vin2 Comparator_0/AND3IN_0/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1071 Comparator_0/OR4IN_0/vin2 Comparator_0/AND3IN_0/NOT_0/in vdd Comparator_0/AND3IN_0/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1072 Comparator_0/AND3IN_0/NOT_0/in Enable_1/vouta2 vdd Comparator_0/AND3IN_0/w_n14_n10# CMOSP w=4 l=2
+  ad=60 pd=54 as=0 ps=0
M1073 Comparator_0/AND3IN_0/a_19_n30# Comparator_0/NOT_1/out Comparator_0/AND3IN_0/a_2_n30# Gnd CMOSN w=4 l=2
+  ad=60 pd=38 as=60 ps=38
M1074 Comparator_0/AND3IN_0/NOT_0/in Comparator_0/NOT_1/out vdd Comparator_0/AND3IN_0/w_n14_n10# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1075 Comparator_0/AND3IN_0/NOT_0/in Comparator_0/NOT_5/out Comparator_0/AND3IN_0/a_19_n30# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1076 Comparator_0/AND3IN_0/a_2_n30# Enable_1/vouta2 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1077 Comparator_0/AND3IN_0/NOT_0/in Comparator_0/NOT_5/out vdd Comparator_0/AND3IN_0/w_n14_n10# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1078 Comparator_0/XOR2IN_0/NAND2IN_0/a_n1_n23# Enable_1/vouta0 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1079 Comparator_0/XOR2IN_0/NAND2IN_2/vin2 Enable_1/vouta0 vdd Comparator_0/XOR2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1080 Comparator_0/XOR2IN_0/NAND2IN_2/vin2 Enable_1/voutb0 Comparator_0/XOR2IN_0/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1081 Comparator_0/XOR2IN_0/NAND2IN_2/vin2 Enable_1/voutb0 vdd Comparator_0/XOR2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1082 Comparator_0/XOR2IN_0/NAND2IN_1/a_n1_n23# Enable_1/vouta0 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1083 Comparator_0/XOR2IN_0/NAND2IN_3/vin1 Enable_1/vouta0 vdd Comparator_0/XOR2IN_0/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1084 Comparator_0/XOR2IN_0/NAND2IN_3/vin1 Comparator_0/XOR2IN_0/NAND2IN_2/vin2 Comparator_0/XOR2IN_0/NAND2IN_1/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1085 Comparator_0/XOR2IN_0/NAND2IN_3/vin1 Comparator_0/XOR2IN_0/NAND2IN_2/vin2 vdd Comparator_0/XOR2IN_0/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1086 Comparator_0/XOR2IN_0/NAND2IN_2/a_n1_n23# Enable_1/voutb0 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1087 Comparator_0/XOR2IN_0/NAND2IN_3/vin2 Enable_1/voutb0 vdd Comparator_0/XOR2IN_0/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1088 Comparator_0/XOR2IN_0/NAND2IN_3/vin2 Comparator_0/XOR2IN_0/NAND2IN_2/vin2 Comparator_0/XOR2IN_0/NAND2IN_2/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1089 Comparator_0/XOR2IN_0/NAND2IN_3/vin2 Comparator_0/XOR2IN_0/NAND2IN_2/vin2 vdd Comparator_0/XOR2IN_0/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1090 Comparator_0/XOR2IN_0/NAND2IN_3/a_n1_n23# Comparator_0/XOR2IN_0/NAND2IN_3/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1091 Comparator_0/NOT_7/in Comparator_0/XOR2IN_0/NAND2IN_3/vin1 vdd Comparator_0/XOR2IN_0/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1092 Comparator_0/NOT_7/in Comparator_0/XOR2IN_0/NAND2IN_3/vin2 Comparator_0/XOR2IN_0/NAND2IN_3/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1093 Comparator_0/NOT_7/in Comparator_0/XOR2IN_0/NAND2IN_3/vin2 vdd Comparator_0/XOR2IN_0/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1094 Comparator_0/XOR2IN_1/NAND2IN_0/a_n1_n23# Enable_1/vouta1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1095 Comparator_0/XOR2IN_1/NAND2IN_2/vin2 Enable_1/vouta1 vdd Comparator_0/XOR2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1096 Comparator_0/XOR2IN_1/NAND2IN_2/vin2 Enable_1/voutb1 Comparator_0/XOR2IN_1/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1097 Comparator_0/XOR2IN_1/NAND2IN_2/vin2 Enable_1/voutb1 vdd Comparator_0/XOR2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1098 Comparator_0/XOR2IN_1/NAND2IN_1/a_n1_n23# Enable_1/vouta1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1099 Comparator_0/XOR2IN_1/NAND2IN_3/vin1 Enable_1/vouta1 vdd Comparator_0/XOR2IN_1/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1100 Comparator_0/XOR2IN_1/NAND2IN_3/vin1 Comparator_0/XOR2IN_1/NAND2IN_2/vin2 Comparator_0/XOR2IN_1/NAND2IN_1/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1101 Comparator_0/XOR2IN_1/NAND2IN_3/vin1 Comparator_0/XOR2IN_1/NAND2IN_2/vin2 vdd Comparator_0/XOR2IN_1/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1102 Comparator_0/XOR2IN_1/NAND2IN_2/a_n1_n23# Enable_1/voutb1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1103 Comparator_0/XOR2IN_1/NAND2IN_3/vin2 Enable_1/voutb1 vdd Comparator_0/XOR2IN_1/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1104 Comparator_0/XOR2IN_1/NAND2IN_3/vin2 Comparator_0/XOR2IN_1/NAND2IN_2/vin2 Comparator_0/XOR2IN_1/NAND2IN_2/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1105 Comparator_0/XOR2IN_1/NAND2IN_3/vin2 Comparator_0/XOR2IN_1/NAND2IN_2/vin2 vdd Comparator_0/XOR2IN_1/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1106 Comparator_0/XOR2IN_1/NAND2IN_3/a_n1_n23# Comparator_0/XOR2IN_1/NAND2IN_3/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1107 Comparator_0/NOT_6/in Comparator_0/XOR2IN_1/NAND2IN_3/vin1 vdd Comparator_0/XOR2IN_1/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1108 Comparator_0/NOT_6/in Comparator_0/XOR2IN_1/NAND2IN_3/vin2 Comparator_0/XOR2IN_1/NAND2IN_3/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1109 Comparator_0/NOT_6/in Comparator_0/XOR2IN_1/NAND2IN_3/vin2 vdd Comparator_0/XOR2IN_1/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1110 Comparator_0/XOR2IN_2/NAND2IN_0/a_n1_n23# Enable_1/vouta2 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1111 Comparator_0/XOR2IN_2/NAND2IN_2/vin2 Enable_1/vouta2 vdd Comparator_0/XOR2IN_2/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1112 Comparator_0/XOR2IN_2/NAND2IN_2/vin2 Enable_1/voutb2 Comparator_0/XOR2IN_2/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1113 Comparator_0/XOR2IN_2/NAND2IN_2/vin2 Enable_1/voutb2 vdd Comparator_0/XOR2IN_2/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1114 Comparator_0/XOR2IN_2/NAND2IN_1/a_n1_n23# Enable_1/vouta2 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1115 Comparator_0/XOR2IN_2/NAND2IN_3/vin1 Enable_1/vouta2 vdd Comparator_0/XOR2IN_2/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1116 Comparator_0/XOR2IN_2/NAND2IN_3/vin1 Comparator_0/XOR2IN_2/NAND2IN_2/vin2 Comparator_0/XOR2IN_2/NAND2IN_1/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1117 Comparator_0/XOR2IN_2/NAND2IN_3/vin1 Comparator_0/XOR2IN_2/NAND2IN_2/vin2 vdd Comparator_0/XOR2IN_2/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1118 Comparator_0/XOR2IN_2/NAND2IN_2/a_n1_n23# Enable_1/voutb2 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1119 Comparator_0/XOR2IN_2/NAND2IN_3/vin2 Enable_1/voutb2 vdd Comparator_0/XOR2IN_2/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1120 Comparator_0/XOR2IN_2/NAND2IN_3/vin2 Comparator_0/XOR2IN_2/NAND2IN_2/vin2 Comparator_0/XOR2IN_2/NAND2IN_2/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1121 Comparator_0/XOR2IN_2/NAND2IN_3/vin2 Comparator_0/XOR2IN_2/NAND2IN_2/vin2 vdd Comparator_0/XOR2IN_2/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1122 Comparator_0/XOR2IN_2/NAND2IN_3/a_n1_n23# Comparator_0/XOR2IN_2/NAND2IN_3/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1123 Comparator_0/NOT_4/in Comparator_0/XOR2IN_2/NAND2IN_3/vin1 vdd Comparator_0/XOR2IN_2/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1124 Comparator_0/NOT_4/in Comparator_0/XOR2IN_2/NAND2IN_3/vin2 Comparator_0/XOR2IN_2/NAND2IN_3/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1125 Comparator_0/NOT_4/in Comparator_0/XOR2IN_2/NAND2IN_3/vin2 vdd Comparator_0/XOR2IN_2/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1126 Comparator_0/XOR2IN_3/NAND2IN_0/a_n1_n23# Enable_1/vouta3 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1127 Comparator_0/XOR2IN_3/NAND2IN_2/vin2 Enable_1/vouta3 vdd Comparator_0/XOR2IN_3/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1128 Comparator_0/XOR2IN_3/NAND2IN_2/vin2 Enable_1/voutb3 Comparator_0/XOR2IN_3/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1129 Comparator_0/XOR2IN_3/NAND2IN_2/vin2 Enable_1/voutb3 vdd Comparator_0/XOR2IN_3/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1130 Comparator_0/XOR2IN_3/NAND2IN_1/a_n1_n23# Enable_1/vouta3 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1131 Comparator_0/XOR2IN_3/NAND2IN_3/vin1 Enable_1/vouta3 vdd Comparator_0/XOR2IN_3/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1132 Comparator_0/XOR2IN_3/NAND2IN_3/vin1 Comparator_0/XOR2IN_3/NAND2IN_2/vin2 Comparator_0/XOR2IN_3/NAND2IN_1/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1133 Comparator_0/XOR2IN_3/NAND2IN_3/vin1 Comparator_0/XOR2IN_3/NAND2IN_2/vin2 vdd Comparator_0/XOR2IN_3/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1134 Comparator_0/XOR2IN_3/NAND2IN_2/a_n1_n23# Enable_1/voutb3 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1135 Comparator_0/XOR2IN_3/NAND2IN_3/vin2 Enable_1/voutb3 vdd Comparator_0/XOR2IN_3/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1136 Comparator_0/XOR2IN_3/NAND2IN_3/vin2 Comparator_0/XOR2IN_3/NAND2IN_2/vin2 Comparator_0/XOR2IN_3/NAND2IN_2/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1137 Comparator_0/XOR2IN_3/NAND2IN_3/vin2 Comparator_0/XOR2IN_3/NAND2IN_2/vin2 vdd Comparator_0/XOR2IN_3/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1138 Comparator_0/XOR2IN_3/NAND2IN_3/a_n1_n23# Comparator_0/XOR2IN_3/NAND2IN_3/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1139 Comparator_0/NOT_5/in Comparator_0/XOR2IN_3/NAND2IN_3/vin1 vdd Comparator_0/XOR2IN_3/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1140 Comparator_0/NOT_5/in Comparator_0/XOR2IN_3/NAND2IN_3/vin2 Comparator_0/XOR2IN_3/NAND2IN_3/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1141 Comparator_0/NOT_5/in Comparator_0/XOR2IN_3/NAND2IN_3/vin2 vdd Comparator_0/XOR2IN_3/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1142 Comparator_0/NOR2IN_0/vout OR3IN_2/vin2 Comparator_0/NOR2IN_0/a_0_1# Comparator_0/NOR2IN_0/w_n19_n9# CMOSP w=12 l=2
+  ad=72 pd=36 as=48 ps=32
M1143 Comparator_0/NOR2IN_0/vout OR3IN_2/vin2 gnd Gnd CMOSN w=4 l=2
+  ad=60 pd=46 as=0 ps=0
M1144 Comparator_0/NOR2IN_0/a_0_1# OR3IN_0/vin2 vdd Comparator_0/NOR2IN_0/w_n19_n9# CMOSP w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1145 Comparator_0/NOR2IN_0/vout OR3IN_0/vin2 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1146 Comparator_0/AND2IN_0/NAND2IN_0/a_n1_n23# Enable_1/vouta3 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1147 Comparator_0/AND2IN_0/NOT_0/in Enable_1/vouta3 vdd Comparator_0/AND2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1148 Comparator_0/AND2IN_0/NOT_0/in Comparator_0/NOT_0/out Comparator_0/AND2IN_0/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1149 Comparator_0/AND2IN_0/NOT_0/in Comparator_0/NOT_0/out vdd Comparator_0/AND2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1150 Comparator_0/OR4IN_0/vin1 Comparator_0/AND2IN_0/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1151 Comparator_0/OR4IN_0/vin1 Comparator_0/AND2IN_0/NOT_0/in vdd Comparator_0/AND2IN_0/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1152 Comparator_0/AND2IN_1/NAND2IN_0/a_n1_n23# Enable_1/vinEn gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1153 Comparator_0/AND2IN_1/NOT_0/in Enable_1/vinEn vdd Comparator_0/AND2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1154 Comparator_0/AND2IN_1/NOT_0/in Comparator_0/AND4IN_0/vout Comparator_0/AND2IN_1/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1155 Comparator_0/AND2IN_1/NOT_0/in Comparator_0/AND4IN_0/vout vdd Comparator_0/AND2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1156 OR3IN_0/vin2 Comparator_0/AND2IN_1/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1157 OR3IN_0/vin2 Comparator_0/AND2IN_1/NOT_0/in vdd Comparator_0/AND2IN_1/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1158 Comparator_0/AND2IN_2/NAND2IN_0/a_n1_n23# Enable_1/vinEn gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1159 Comparator_0/AND2IN_2/NOT_0/in Enable_1/vinEn vdd Comparator_0/AND2IN_2/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1160 Comparator_0/AND2IN_2/NOT_0/in Comparator_0/OR4IN_0/vout Comparator_0/AND2IN_2/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1161 Comparator_0/AND2IN_2/NOT_0/in Comparator_0/OR4IN_0/vout vdd Comparator_0/AND2IN_2/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1162 OR3IN_2/vin2 Comparator_0/AND2IN_2/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1163 OR3IN_2/vin2 Comparator_0/AND2IN_2/NOT_0/in vdd Comparator_0/AND2IN_2/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=55 pd=42 as=0 ps=0
M1164 Comparator_0/OR4IN_0/vin4 Comparator_0/AND5IN_0/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1165 Comparator_0/OR4IN_0/vin4 Comparator_0/AND5IN_0/NOT_0/in vdd Comparator_0/AND5IN_0/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1166 Comparator_0/AND5IN_0/NOT_0/in Comparator_0/NOT_5/out vdd Comparator_0/AND5IN_0/w_n26_1# CMOSP w=4 l=2
+  ad=100 pd=90 as=0 ps=0
M1167 Comparator_0/AND5IN_0/NOT_0/in Comparator_0/NOT_6/out Comparator_0/AND5IN_0/a_36_n32# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=56 ps=36
M1168 Comparator_0/AND5IN_0/a_20_n32# Comparator_0/NOT_5/out Comparator_0/AND5IN_0/a_4_n32# Gnd CMOSN w=4 l=2
+  ad=56 pd=36 as=56 ps=36
M1169 Comparator_0/AND5IN_0/NOT_0/in Comparator_0/NOT_3/out vdd Comparator_0/AND5IN_0/w_n26_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1170 Comparator_0/AND5IN_0/a_4_n32# Comparator_0/NOT_3/out Comparator_0/AND5IN_0/a_n12_n32# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=56 ps=36
M1171 Comparator_0/AND5IN_0/NOT_0/in Comparator_0/NOT_6/out vdd Comparator_0/AND5IN_0/w_n26_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1172 Comparator_0/AND5IN_0/a_n12_n32# Enable_1/vouta0 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1173 Comparator_0/AND5IN_0/NOT_0/in Enable_1/vouta0 vdd Comparator_0/AND5IN_0/w_n26_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1174 Comparator_0/AND5IN_0/a_36_n32# Comparator_0/NOT_4/out Comparator_0/AND5IN_0/a_20_n32# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1175 Comparator_0/AND5IN_0/NOT_0/in Comparator_0/NOT_4/out vdd Comparator_0/AND5IN_0/w_n26_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1176 Comparator_0/AND2IN_3/NAND2IN_0/a_n1_n23# Comparator_0/NOR2IN_0/vout gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1177 Comparator_0/AND2IN_3/NOT_0/in Comparator_0/NOR2IN_0/vout vdd Comparator_0/AND2IN_3/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1178 Comparator_0/AND2IN_3/NOT_0/in Enable_1/vinEn Comparator_0/AND2IN_3/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1179 Comparator_0/AND2IN_3/NOT_0/in Enable_1/vinEn vdd Comparator_0/AND2IN_3/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1180 OR3IN_1/vin2 Comparator_0/AND2IN_3/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1181 OR3IN_1/vin2 Comparator_0/AND2IN_3/NOT_0/in vdd Comparator_0/AND2IN_3/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1182 Comparator_0/NOT_1/out Enable_1/voutb2 gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1183 Comparator_0/NOT_1/out Enable_1/voutb2 vdd Comparator_0/NOT_1/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1184 Comparator_0/NOT_0/out Enable_1/voutb3 gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1185 Comparator_0/NOT_0/out Enable_1/voutb3 vdd Comparator_0/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1186 Comparator_0/NOT_2/out Enable_1/voutb1 gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1187 Comparator_0/NOT_2/out Enable_1/voutb1 vdd Comparator_0/NOT_2/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1188 Comparator_0/AND4IN_0/vout Comparator_0/AND4IN_0/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1189 Comparator_0/AND4IN_0/vout Comparator_0/AND4IN_0/NOT_0/in vdd Comparator_0/AND4IN_0/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1190 Comparator_0/AND4IN_0/NOT_0/in Comparator_0/NOT_7/out vdd Comparator_0/AND4IN_0/w_n14_n10# CMOSP w=4 l=2
+  ad=80 pd=72 as=0 ps=0
M1191 Comparator_0/AND4IN_0/a_19_n30# Comparator_0/NOT_6/out Comparator_0/AND4IN_0/a_2_n30# Gnd CMOSN w=4 l=2
+  ad=60 pd=38 as=60 ps=38
M1192 Comparator_0/AND4IN_0/NOT_0/in Comparator_0/NOT_5/out vdd Comparator_0/AND4IN_0/w_n14_n10# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1193 Comparator_0/AND4IN_0/NOT_0/in Comparator_0/NOT_6/out vdd Comparator_0/AND4IN_0/w_n14_n10# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1194 Comparator_0/AND4IN_0/a_36_n30# Comparator_0/NOT_4/out Comparator_0/AND4IN_0/a_19_n30# Gnd CMOSN w=4 l=2
+  ad=60 pd=38 as=0 ps=0
M1195 Comparator_0/AND4IN_0/NOT_0/in Comparator_0/NOT_5/out Comparator_0/AND4IN_0/a_36_n30# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1196 Comparator_0/AND4IN_0/a_2_n30# Comparator_0/NOT_7/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1197 Comparator_0/AND4IN_0/NOT_0/in Comparator_0/NOT_4/out vdd Comparator_0/AND4IN_0/w_n14_n10# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1198 Comparator_0/NOT_3/out Enable_1/voutb0 gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1199 Comparator_0/NOT_3/out Enable_1/voutb0 vdd Comparator_0/NOT_3/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1200 Comparator_0/OR4IN_0/vin3 Comparator_0/AND4IN_1/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1201 Comparator_0/OR4IN_0/vin3 Comparator_0/AND4IN_1/NOT_0/in vdd Comparator_0/AND4IN_1/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1202 Comparator_0/AND4IN_1/NOT_0/in Enable_1/vouta1 vdd Comparator_0/AND4IN_1/w_n14_n10# CMOSP w=4 l=2
+  ad=80 pd=72 as=0 ps=0
M1203 Comparator_0/AND4IN_1/a_19_n30# Comparator_0/NOT_2/out Comparator_0/AND4IN_1/a_2_n30# Gnd CMOSN w=4 l=2
+  ad=60 pd=38 as=60 ps=38
M1204 Comparator_0/AND4IN_1/NOT_0/in Comparator_0/NOT_4/out vdd Comparator_0/AND4IN_1/w_n14_n10# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1205 Comparator_0/AND4IN_1/NOT_0/in Comparator_0/NOT_2/out vdd Comparator_0/AND4IN_1/w_n14_n10# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1206 Comparator_0/AND4IN_1/a_36_n30# Comparator_0/NOT_5/out Comparator_0/AND4IN_1/a_19_n30# Gnd CMOSN w=4 l=2
+  ad=60 pd=38 as=0 ps=0
M1207 Comparator_0/AND4IN_1/NOT_0/in Comparator_0/NOT_4/out Comparator_0/AND4IN_1/a_36_n30# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1208 Comparator_0/AND4IN_1/a_2_n30# Enable_1/vouta1 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1209 Comparator_0/AND4IN_1/NOT_0/in Comparator_0/NOT_5/out vdd Comparator_0/AND4IN_1/w_n14_n10# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1210 Comparator_0/NOT_4/out Comparator_0/NOT_4/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1211 Comparator_0/NOT_4/out Comparator_0/NOT_4/in vdd Comparator_0/NOT_4/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1212 Comparator_0/OR4IN_0/vout Comparator_0/OR4IN_0/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1213 Comparator_0/OR4IN_0/vout Comparator_0/OR4IN_0/NOT_0/in vdd Comparator_0/OR4IN_0/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1214 Comparator_0/OR4IN_0/a_6_1# Comparator_0/OR4IN_0/vin2 Comparator_0/OR4IN_0/a_0_1# Comparator_0/OR4IN_0/w_n19_n9# CMOSP w=12 l=2
+  ad=48 pd=32 as=48 ps=32
M1215 Comparator_0/OR4IN_0/a_0_1# Comparator_0/OR4IN_0/vin1 vdd Comparator_0/OR4IN_0/w_n19_n9# CMOSP w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1216 Comparator_0/OR4IN_0/NOT_0/in Comparator_0/OR4IN_0/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=112 pd=88 as=0 ps=0
M1217 Comparator_0/OR4IN_0/NOT_0/in Comparator_0/OR4IN_0/vin3 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1218 Comparator_0/OR4IN_0/NOT_0/in Comparator_0/OR4IN_0/vin4 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1219 Comparator_0/OR4IN_0/NOT_0/in Comparator_0/OR4IN_0/vin4 Comparator_0/OR4IN_0/a_12_1# Comparator_0/OR4IN_0/w_n19_n9# CMOSP w=12 l=2
+  ad=120 pd=44 as=48 ps=32
M1220 Comparator_0/OR4IN_0/a_12_1# Comparator_0/OR4IN_0/vin3 Comparator_0/OR4IN_0/a_6_1# Comparator_0/OR4IN_0/w_n19_n9# CMOSP w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1221 Comparator_0/OR4IN_0/NOT_0/in Comparator_0/OR4IN_0/vin2 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1222 AND4Bit_0/AND2IN_0/NAND2IN_0/a_n1_n23# Enable_2/vouta0 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1223 AND4Bit_0/AND2IN_0/NOT_0/in Enable_2/vouta0 vdd AND4Bit_0/AND2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1224 AND4Bit_0/AND2IN_0/NOT_0/in Enable_2/voutb0 AND4Bit_0/AND2IN_0/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1225 AND4Bit_0/AND2IN_0/NOT_0/in Enable_2/voutb0 vdd AND4Bit_0/AND2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1226 OR3IN_0/vin3 AND4Bit_0/AND2IN_0/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1227 OR3IN_0/vin3 AND4Bit_0/AND2IN_0/NOT_0/in vdd AND4Bit_0/AND2IN_0/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1228 AND4Bit_0/AND2IN_1/NAND2IN_0/a_n1_n23# Enable_2/vouta1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1229 AND4Bit_0/AND2IN_1/NOT_0/in Enable_2/vouta1 vdd AND4Bit_0/AND2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1230 AND4Bit_0/AND2IN_1/NOT_0/in Enable_2/voutb1 AND4Bit_0/AND2IN_1/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1231 AND4Bit_0/AND2IN_1/NOT_0/in Enable_2/voutb1 vdd AND4Bit_0/AND2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1232 OR3IN_1/vin3 AND4Bit_0/AND2IN_1/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1233 OR3IN_1/vin3 AND4Bit_0/AND2IN_1/NOT_0/in vdd AND4Bit_0/AND2IN_1/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1234 AND4Bit_0/AND2IN_2/NAND2IN_0/a_n1_n23# Enable_2/vouta2 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1235 AND4Bit_0/AND2IN_2/NOT_0/in Enable_2/vouta2 vdd AND4Bit_0/AND2IN_2/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1236 AND4Bit_0/AND2IN_2/NOT_0/in Enable_2/voutb2 AND4Bit_0/AND2IN_2/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1237 AND4Bit_0/AND2IN_2/NOT_0/in Enable_2/voutb2 vdd AND4Bit_0/AND2IN_2/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1238 OR3IN_2/vin3 AND4Bit_0/AND2IN_2/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1239 OR3IN_2/vin3 AND4Bit_0/AND2IN_2/NOT_0/in vdd AND4Bit_0/AND2IN_2/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1240 AND4Bit_0/AND2IN_3/NAND2IN_0/a_n1_n23# Enable_2/vouta3 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1241 AND4Bit_0/AND2IN_3/NOT_0/in Enable_2/vouta3 vdd AND4Bit_0/AND2IN_3/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1242 AND4Bit_0/AND2IN_3/NOT_0/in Enable_2/voutb3 AND4Bit_0/AND2IN_3/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1243 AND4Bit_0/AND2IN_3/NOT_0/in Enable_2/voutb3 vdd AND4Bit_0/AND2IN_3/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1244 OR2IN_1/vin2 AND4Bit_0/AND2IN_3/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1245 OR2IN_1/vin2 AND4Bit_0/AND2IN_3/NOT_0/in vdd AND4Bit_0/AND2IN_3/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1246 Enable_0/AND4Bit_0/AND2IN_0/NAND2IN_0/a_n1_n23# vina0 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1247 Enable_0/AND4Bit_0/AND2IN_0/NOT_0/in vina0 vdd Enable_0/AND4Bit_0/AND2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1248 Enable_0/AND4Bit_0/AND2IN_0/NOT_0/in OR2IN_0/vout Enable_0/AND4Bit_0/AND2IN_0/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1249 Enable_0/AND4Bit_0/AND2IN_0/NOT_0/in OR2IN_0/vout vdd Enable_0/AND4Bit_0/AND2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1250 Enable_0/vouta0 Enable_0/AND4Bit_0/AND2IN_0/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1251 Enable_0/vouta0 Enable_0/AND4Bit_0/AND2IN_0/NOT_0/in vdd Enable_0/AND4Bit_0/AND2IN_0/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1252 Enable_0/AND4Bit_0/AND2IN_1/NAND2IN_0/a_n1_n23# vina1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1253 Enable_0/AND4Bit_0/AND2IN_1/NOT_0/in vina1 vdd Enable_0/AND4Bit_0/AND2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1254 Enable_0/AND4Bit_0/AND2IN_1/NOT_0/in OR2IN_0/vout Enable_0/AND4Bit_0/AND2IN_1/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1255 Enable_0/AND4Bit_0/AND2IN_1/NOT_0/in OR2IN_0/vout vdd Enable_0/AND4Bit_0/AND2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1256 Enable_0/vouta1 Enable_0/AND4Bit_0/AND2IN_1/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1257 Enable_0/vouta1 Enable_0/AND4Bit_0/AND2IN_1/NOT_0/in vdd Enable_0/AND4Bit_0/AND2IN_1/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1258 Enable_0/AND4Bit_0/AND2IN_2/NAND2IN_0/a_n1_n23# vina2 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1259 Enable_0/AND4Bit_0/AND2IN_2/NOT_0/in vina2 vdd Enable_0/AND4Bit_0/AND2IN_2/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1260 Enable_0/AND4Bit_0/AND2IN_2/NOT_0/in OR2IN_0/vout Enable_0/AND4Bit_0/AND2IN_2/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1261 Enable_0/AND4Bit_0/AND2IN_2/NOT_0/in OR2IN_0/vout vdd Enable_0/AND4Bit_0/AND2IN_2/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1262 Enable_0/vouta2 Enable_0/AND4Bit_0/AND2IN_2/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1263 Enable_0/vouta2 Enable_0/AND4Bit_0/AND2IN_2/NOT_0/in vdd Enable_0/AND4Bit_0/AND2IN_2/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1264 Enable_0/AND4Bit_0/AND2IN_3/NAND2IN_0/a_n1_n23# vina3 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1265 Enable_0/AND4Bit_0/AND2IN_3/NOT_0/in vina3 vdd Enable_0/AND4Bit_0/AND2IN_3/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1266 Enable_0/AND4Bit_0/AND2IN_3/NOT_0/in OR2IN_0/vout Enable_0/AND4Bit_0/AND2IN_3/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1267 Enable_0/AND4Bit_0/AND2IN_3/NOT_0/in OR2IN_0/vout vdd Enable_0/AND4Bit_0/AND2IN_3/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1268 Enable_0/vouta3 Enable_0/AND4Bit_0/AND2IN_3/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1269 Enable_0/vouta3 Enable_0/AND4Bit_0/AND2IN_3/NOT_0/in vdd Enable_0/AND4Bit_0/AND2IN_3/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1270 Enable_0/AND4Bit_1/AND2IN_0/NAND2IN_0/a_n1_n23# vinb0 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1271 Enable_0/AND4Bit_1/AND2IN_0/NOT_0/in vinb0 vdd Enable_0/AND4Bit_1/AND2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1272 Enable_0/AND4Bit_1/AND2IN_0/NOT_0/in OR2IN_0/vout Enable_0/AND4Bit_1/AND2IN_0/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1273 Enable_0/AND4Bit_1/AND2IN_0/NOT_0/in OR2IN_0/vout vdd Enable_0/AND4Bit_1/AND2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1274 Enable_0/voutb0 Enable_0/AND4Bit_1/AND2IN_0/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1275 Enable_0/voutb0 Enable_0/AND4Bit_1/AND2IN_0/NOT_0/in vdd Enable_0/AND4Bit_1/AND2IN_0/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1276 Enable_0/AND4Bit_1/AND2IN_1/NAND2IN_0/a_n1_n23# vinb1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1277 Enable_0/AND4Bit_1/AND2IN_1/NOT_0/in vinb1 vdd Enable_0/AND4Bit_1/AND2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1278 Enable_0/AND4Bit_1/AND2IN_1/NOT_0/in OR2IN_0/vout Enable_0/AND4Bit_1/AND2IN_1/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1279 Enable_0/AND4Bit_1/AND2IN_1/NOT_0/in OR2IN_0/vout vdd Enable_0/AND4Bit_1/AND2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1280 Enable_0/voutb1 Enable_0/AND4Bit_1/AND2IN_1/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1281 Enable_0/voutb1 Enable_0/AND4Bit_1/AND2IN_1/NOT_0/in vdd Enable_0/AND4Bit_1/AND2IN_1/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1282 Enable_0/AND4Bit_1/AND2IN_2/NAND2IN_0/a_n1_n23# vinb2 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1283 Enable_0/AND4Bit_1/AND2IN_2/NOT_0/in vinb2 vdd Enable_0/AND4Bit_1/AND2IN_2/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1284 Enable_0/AND4Bit_1/AND2IN_2/NOT_0/in OR2IN_0/vout Enable_0/AND4Bit_1/AND2IN_2/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1285 Enable_0/AND4Bit_1/AND2IN_2/NOT_0/in OR2IN_0/vout vdd Enable_0/AND4Bit_1/AND2IN_2/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1286 Enable_0/voutb2 Enable_0/AND4Bit_1/AND2IN_2/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1287 Enable_0/voutb2 Enable_0/AND4Bit_1/AND2IN_2/NOT_0/in vdd Enable_0/AND4Bit_1/AND2IN_2/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1288 Enable_0/AND4Bit_1/AND2IN_3/NAND2IN_0/a_n1_n23# vinb3 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1289 Enable_0/AND4Bit_1/AND2IN_3/NOT_0/in vinb3 vdd Enable_0/AND4Bit_1/AND2IN_3/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1290 Enable_0/AND4Bit_1/AND2IN_3/NOT_0/in OR2IN_0/vout Enable_0/AND4Bit_1/AND2IN_3/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1291 Enable_0/AND4Bit_1/AND2IN_3/NOT_0/in OR2IN_0/vout vdd Enable_0/AND4Bit_1/AND2IN_3/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1292 Enable_0/voutb3 Enable_0/AND4Bit_1/AND2IN_3/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1293 Enable_0/voutb3 Enable_0/AND4Bit_1/AND2IN_3/NOT_0/in vdd Enable_0/AND4Bit_1/AND2IN_3/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1294 Enable_1/AND4Bit_0/AND2IN_0/NAND2IN_0/a_n1_n23# vina0 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1295 Enable_1/AND4Bit_0/AND2IN_0/NOT_0/in vina0 vdd Enable_1/AND4Bit_0/AND2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1296 Enable_1/AND4Bit_0/AND2IN_0/NOT_0/in Enable_1/vinEn Enable_1/AND4Bit_0/AND2IN_0/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1297 Enable_1/AND4Bit_0/AND2IN_0/NOT_0/in Enable_1/vinEn vdd Enable_1/AND4Bit_0/AND2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1298 Enable_1/vouta0 Enable_1/AND4Bit_0/AND2IN_0/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1299 Enable_1/vouta0 Enable_1/AND4Bit_0/AND2IN_0/NOT_0/in vdd Enable_1/AND4Bit_0/AND2IN_0/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1300 Enable_1/AND4Bit_0/AND2IN_1/NAND2IN_0/a_n1_n23# vina1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1301 Enable_1/AND4Bit_0/AND2IN_1/NOT_0/in vina1 vdd Enable_1/AND4Bit_0/AND2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1302 Enable_1/AND4Bit_0/AND2IN_1/NOT_0/in Enable_1/vinEn Enable_1/AND4Bit_0/AND2IN_1/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1303 Enable_1/AND4Bit_0/AND2IN_1/NOT_0/in Enable_1/vinEn vdd Enable_1/AND4Bit_0/AND2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1304 Enable_1/vouta1 Enable_1/AND4Bit_0/AND2IN_1/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1305 Enable_1/vouta1 Enable_1/AND4Bit_0/AND2IN_1/NOT_0/in vdd Enable_1/AND4Bit_0/AND2IN_1/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1306 Enable_1/AND4Bit_0/AND2IN_2/NAND2IN_0/a_n1_n23# vina2 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1307 Enable_1/AND4Bit_0/AND2IN_2/NOT_0/in vina2 vdd Enable_1/AND4Bit_0/AND2IN_2/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1308 Enable_1/AND4Bit_0/AND2IN_2/NOT_0/in Enable_1/vinEn Enable_1/AND4Bit_0/AND2IN_2/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1309 Enable_1/AND4Bit_0/AND2IN_2/NOT_0/in Enable_1/vinEn vdd Enable_1/AND4Bit_0/AND2IN_2/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1310 Enable_1/vouta2 Enable_1/AND4Bit_0/AND2IN_2/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1311 Enable_1/vouta2 Enable_1/AND4Bit_0/AND2IN_2/NOT_0/in vdd Enable_1/AND4Bit_0/AND2IN_2/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1312 Enable_1/AND4Bit_0/AND2IN_3/NAND2IN_0/a_n1_n23# vina3 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1313 Enable_1/AND4Bit_0/AND2IN_3/NOT_0/in vina3 vdd Enable_1/AND4Bit_0/AND2IN_3/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1314 Enable_1/AND4Bit_0/AND2IN_3/NOT_0/in Enable_1/vinEn Enable_1/AND4Bit_0/AND2IN_3/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1315 Enable_1/AND4Bit_0/AND2IN_3/NOT_0/in Enable_1/vinEn vdd Enable_1/AND4Bit_0/AND2IN_3/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1316 Enable_1/vouta3 Enable_1/AND4Bit_0/AND2IN_3/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1317 Enable_1/vouta3 Enable_1/AND4Bit_0/AND2IN_3/NOT_0/in vdd Enable_1/AND4Bit_0/AND2IN_3/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1318 Enable_1/AND4Bit_1/AND2IN_0/NAND2IN_0/a_n1_n23# vinb0 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1319 Enable_1/AND4Bit_1/AND2IN_0/NOT_0/in vinb0 vdd Enable_1/AND4Bit_1/AND2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1320 Enable_1/AND4Bit_1/AND2IN_0/NOT_0/in Enable_1/vinEn Enable_1/AND4Bit_1/AND2IN_0/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1321 Enable_1/AND4Bit_1/AND2IN_0/NOT_0/in Enable_1/vinEn vdd Enable_1/AND4Bit_1/AND2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1322 Enable_1/voutb0 Enable_1/AND4Bit_1/AND2IN_0/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1323 Enable_1/voutb0 Enable_1/AND4Bit_1/AND2IN_0/NOT_0/in vdd Enable_1/AND4Bit_1/AND2IN_0/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1324 Enable_1/AND4Bit_1/AND2IN_1/NAND2IN_0/a_n1_n23# vinb1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1325 Enable_1/AND4Bit_1/AND2IN_1/NOT_0/in vinb1 vdd Enable_1/AND4Bit_1/AND2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1326 Enable_1/AND4Bit_1/AND2IN_1/NOT_0/in Enable_1/vinEn Enable_1/AND4Bit_1/AND2IN_1/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1327 Enable_1/AND4Bit_1/AND2IN_1/NOT_0/in Enable_1/vinEn vdd Enable_1/AND4Bit_1/AND2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1328 Enable_1/voutb1 Enable_1/AND4Bit_1/AND2IN_1/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1329 Enable_1/voutb1 Enable_1/AND4Bit_1/AND2IN_1/NOT_0/in vdd Enable_1/AND4Bit_1/AND2IN_1/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1330 Enable_1/AND4Bit_1/AND2IN_2/NAND2IN_0/a_n1_n23# vinb2 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1331 Enable_1/AND4Bit_1/AND2IN_2/NOT_0/in vinb2 vdd Enable_1/AND4Bit_1/AND2IN_2/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1332 Enable_1/AND4Bit_1/AND2IN_2/NOT_0/in Enable_1/vinEn Enable_1/AND4Bit_1/AND2IN_2/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1333 Enable_1/AND4Bit_1/AND2IN_2/NOT_0/in Enable_1/vinEn vdd Enable_1/AND4Bit_1/AND2IN_2/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1334 Enable_1/voutb2 Enable_1/AND4Bit_1/AND2IN_2/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1335 Enable_1/voutb2 Enable_1/AND4Bit_1/AND2IN_2/NOT_0/in vdd Enable_1/AND4Bit_1/AND2IN_2/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1336 Enable_1/AND4Bit_1/AND2IN_3/NAND2IN_0/a_n1_n23# vinb3 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1337 Enable_1/AND4Bit_1/AND2IN_3/NOT_0/in vinb3 vdd Enable_1/AND4Bit_1/AND2IN_3/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1338 Enable_1/AND4Bit_1/AND2IN_3/NOT_0/in Enable_1/vinEn Enable_1/AND4Bit_1/AND2IN_3/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1339 Enable_1/AND4Bit_1/AND2IN_3/NOT_0/in Enable_1/vinEn vdd Enable_1/AND4Bit_1/AND2IN_3/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1340 Enable_1/voutb3 Enable_1/AND4Bit_1/AND2IN_3/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1341 Enable_1/voutb3 Enable_1/AND4Bit_1/AND2IN_3/NOT_0/in vdd Enable_1/AND4Bit_1/AND2IN_3/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1342 Enable_2/AND4Bit_0/AND2IN_0/NAND2IN_0/a_n1_n23# vina0 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1343 Enable_2/AND4Bit_0/AND2IN_0/NOT_0/in vina0 vdd Enable_2/AND4Bit_0/AND2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1344 Enable_2/AND4Bit_0/AND2IN_0/NOT_0/in Enable_2/vinEn Enable_2/AND4Bit_0/AND2IN_0/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1345 Enable_2/AND4Bit_0/AND2IN_0/NOT_0/in Enable_2/vinEn vdd Enable_2/AND4Bit_0/AND2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1346 Enable_2/vouta0 Enable_2/AND4Bit_0/AND2IN_0/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1347 Enable_2/vouta0 Enable_2/AND4Bit_0/AND2IN_0/NOT_0/in vdd Enable_2/AND4Bit_0/AND2IN_0/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1348 Enable_2/AND4Bit_0/AND2IN_1/NAND2IN_0/a_n1_n23# vina1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1349 Enable_2/AND4Bit_0/AND2IN_1/NOT_0/in vina1 vdd Enable_2/AND4Bit_0/AND2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1350 Enable_2/AND4Bit_0/AND2IN_1/NOT_0/in Enable_2/vinEn Enable_2/AND4Bit_0/AND2IN_1/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1351 Enable_2/AND4Bit_0/AND2IN_1/NOT_0/in Enable_2/vinEn vdd Enable_2/AND4Bit_0/AND2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1352 Enable_2/vouta1 Enable_2/AND4Bit_0/AND2IN_1/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1353 Enable_2/vouta1 Enable_2/AND4Bit_0/AND2IN_1/NOT_0/in vdd Enable_2/AND4Bit_0/AND2IN_1/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1354 Enable_2/AND4Bit_0/AND2IN_2/NAND2IN_0/a_n1_n23# vina2 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1355 Enable_2/AND4Bit_0/AND2IN_2/NOT_0/in vina2 vdd Enable_2/AND4Bit_0/AND2IN_2/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1356 Enable_2/AND4Bit_0/AND2IN_2/NOT_0/in Enable_2/vinEn Enable_2/AND4Bit_0/AND2IN_2/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1357 Enable_2/AND4Bit_0/AND2IN_2/NOT_0/in Enable_2/vinEn vdd Enable_2/AND4Bit_0/AND2IN_2/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1358 Enable_2/vouta2 Enable_2/AND4Bit_0/AND2IN_2/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1359 Enable_2/vouta2 Enable_2/AND4Bit_0/AND2IN_2/NOT_0/in vdd Enable_2/AND4Bit_0/AND2IN_2/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1360 Enable_2/AND4Bit_0/AND2IN_3/NAND2IN_0/a_n1_n23# vina3 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1361 Enable_2/AND4Bit_0/AND2IN_3/NOT_0/in vina3 vdd Enable_2/AND4Bit_0/AND2IN_3/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1362 Enable_2/AND4Bit_0/AND2IN_3/NOT_0/in Enable_2/vinEn Enable_2/AND4Bit_0/AND2IN_3/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1363 Enable_2/AND4Bit_0/AND2IN_3/NOT_0/in Enable_2/vinEn vdd Enable_2/AND4Bit_0/AND2IN_3/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1364 Enable_2/vouta3 Enable_2/AND4Bit_0/AND2IN_3/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1365 Enable_2/vouta3 Enable_2/AND4Bit_0/AND2IN_3/NOT_0/in vdd Enable_2/AND4Bit_0/AND2IN_3/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1366 Enable_2/AND4Bit_1/AND2IN_0/NAND2IN_0/a_n1_n23# vinb0 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1367 Enable_2/AND4Bit_1/AND2IN_0/NOT_0/in vinb0 vdd Enable_2/AND4Bit_1/AND2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1368 Enable_2/AND4Bit_1/AND2IN_0/NOT_0/in Enable_2/vinEn Enable_2/AND4Bit_1/AND2IN_0/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1369 Enable_2/AND4Bit_1/AND2IN_0/NOT_0/in Enable_2/vinEn vdd Enable_2/AND4Bit_1/AND2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1370 Enable_2/voutb0 Enable_2/AND4Bit_1/AND2IN_0/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1371 Enable_2/voutb0 Enable_2/AND4Bit_1/AND2IN_0/NOT_0/in vdd Enable_2/AND4Bit_1/AND2IN_0/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1372 Enable_2/AND4Bit_1/AND2IN_1/NAND2IN_0/a_n1_n23# vinb1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1373 Enable_2/AND4Bit_1/AND2IN_1/NOT_0/in vinb1 vdd Enable_2/AND4Bit_1/AND2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1374 Enable_2/AND4Bit_1/AND2IN_1/NOT_0/in Enable_2/vinEn Enable_2/AND4Bit_1/AND2IN_1/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1375 Enable_2/AND4Bit_1/AND2IN_1/NOT_0/in Enable_2/vinEn vdd Enable_2/AND4Bit_1/AND2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1376 Enable_2/voutb1 Enable_2/AND4Bit_1/AND2IN_1/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1377 Enable_2/voutb1 Enable_2/AND4Bit_1/AND2IN_1/NOT_0/in vdd Enable_2/AND4Bit_1/AND2IN_1/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1378 Enable_2/AND4Bit_1/AND2IN_2/NAND2IN_0/a_n1_n23# vinb2 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1379 Enable_2/AND4Bit_1/AND2IN_2/NOT_0/in vinb2 vdd Enable_2/AND4Bit_1/AND2IN_2/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1380 Enable_2/AND4Bit_1/AND2IN_2/NOT_0/in Enable_2/vinEn Enable_2/AND4Bit_1/AND2IN_2/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1381 Enable_2/AND4Bit_1/AND2IN_2/NOT_0/in Enable_2/vinEn vdd Enable_2/AND4Bit_1/AND2IN_2/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1382 Enable_2/voutb2 Enable_2/AND4Bit_1/AND2IN_2/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1383 Enable_2/voutb2 Enable_2/AND4Bit_1/AND2IN_2/NOT_0/in vdd Enable_2/AND4Bit_1/AND2IN_2/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1384 Enable_2/AND4Bit_1/AND2IN_3/NAND2IN_0/a_n1_n23# vinb3 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1385 Enable_2/AND4Bit_1/AND2IN_3/NOT_0/in vinb3 vdd Enable_2/AND4Bit_1/AND2IN_3/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1386 Enable_2/AND4Bit_1/AND2IN_3/NOT_0/in Enable_2/vinEn Enable_2/AND4Bit_1/AND2IN_3/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1387 Enable_2/AND4Bit_1/AND2IN_3/NOT_0/in Enable_2/vinEn vdd Enable_2/AND4Bit_1/AND2IN_3/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1388 Enable_2/voutb3 Enable_2/AND4Bit_1/AND2IN_3/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1389 Enable_2/voutb3 Enable_2/AND4Bit_1/AND2IN_3/NOT_0/in vdd Enable_2/AND4Bit_1/AND2IN_3/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1390 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_0/a_n1_n23# AdderSubtractor_0/fullAdder_2/XOR2IN_1/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1391 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_2/XOR2IN_1/vin1 vdd AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1392 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_2/vcin AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1393 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_2/vcin vdd AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1394 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_1/a_n1_n23# AdderSubtractor_0/fullAdder_2/XOR2IN_1/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1395 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_3/vin1 AdderSubtractor_0/fullAdder_2/XOR2IN_1/vin1 vdd AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1396 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_3/vin1 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_1/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1397 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_3/vin1 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_2/vin2 vdd AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1398 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_2/a_n1_n23# AdderSubtractor_0/fullAdder_2/vcin gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1399 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_3/vin2 AdderSubtractor_0/fullAdder_2/vcin vdd AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1400 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_3/vin2 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_2/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1401 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_3/vin2 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_2/vin2 vdd AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1402 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_3/a_n1_n23# AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_3/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1403 OR3IN_2/vin1 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_3/vin1 vdd AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1404 OR3IN_2/vin1 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_3/vin2 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_3/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1405 OR3IN_2/vin1 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_3/vin2 vdd AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1406 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_0/a_n1_n23# Enable_0/vouta2 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1407 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_2/vin2 Enable_0/vouta2 vdd AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1408 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_2/vin2 AdderSubtractor_0/XOR2IN_2/vout AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1409 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_2/vin2 AdderSubtractor_0/XOR2IN_2/vout vdd AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1410 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_1/a_n1_n23# Enable_0/vouta2 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1411 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_3/vin1 Enable_0/vouta2 vdd AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1412 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_3/vin1 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_1/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1413 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_3/vin1 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_2/vin2 vdd AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1414 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_2/a_n1_n23# AdderSubtractor_0/XOR2IN_2/vout gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1415 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_3/vin2 AdderSubtractor_0/XOR2IN_2/vout vdd AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1416 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_3/vin2 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_2/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1417 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_3/vin2 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_2/vin2 vdd AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1418 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_3/a_n1_n23# AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_3/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1419 AdderSubtractor_0/fullAdder_2/XOR2IN_1/vin1 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_3/vin1 vdd AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1420 AdderSubtractor_0/fullAdder_2/XOR2IN_1/vin1 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_3/vin2 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_3/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1421 AdderSubtractor_0/fullAdder_2/XOR2IN_1/vin1 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_3/vin2 vdd AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1422 AdderSubtractor_0/fullAdder_2/AND2IN_0/NAND2IN_0/a_n1_n23# Enable_0/vouta2 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1423 AdderSubtractor_0/fullAdder_2/AND2IN_0/NOT_0/in Enable_0/vouta2 vdd AdderSubtractor_0/fullAdder_2/AND2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1424 AdderSubtractor_0/fullAdder_2/AND2IN_0/NOT_0/in AdderSubtractor_0/XOR2IN_2/vout AdderSubtractor_0/fullAdder_2/AND2IN_0/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1425 AdderSubtractor_0/fullAdder_2/AND2IN_0/NOT_0/in AdderSubtractor_0/XOR2IN_2/vout vdd AdderSubtractor_0/fullAdder_2/AND2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1426 AdderSubtractor_0/fullAdder_2/OR2IN_0/vin2 AdderSubtractor_0/fullAdder_2/AND2IN_0/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1427 AdderSubtractor_0/fullAdder_2/OR2IN_0/vin2 AdderSubtractor_0/fullAdder_2/AND2IN_0/NOT_0/in vdd AdderSubtractor_0/fullAdder_2/AND2IN_0/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1428 AdderSubtractor_0/fullAdder_2/AND2IN_1/NAND2IN_0/a_n1_n23# AdderSubtractor_0/fullAdder_2/vcin gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1429 AdderSubtractor_0/fullAdder_2/AND2IN_1/NOT_0/in AdderSubtractor_0/fullAdder_2/vcin vdd AdderSubtractor_0/fullAdder_2/AND2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1430 AdderSubtractor_0/fullAdder_2/AND2IN_1/NOT_0/in AdderSubtractor_0/fullAdder_2/XOR2IN_1/vin1 AdderSubtractor_0/fullAdder_2/AND2IN_1/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1431 AdderSubtractor_0/fullAdder_2/AND2IN_1/NOT_0/in AdderSubtractor_0/fullAdder_2/XOR2IN_1/vin1 vdd AdderSubtractor_0/fullAdder_2/AND2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1432 AdderSubtractor_0/fullAdder_2/OR2IN_0/vin1 AdderSubtractor_0/fullAdder_2/AND2IN_1/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1433 AdderSubtractor_0/fullAdder_2/OR2IN_0/vin1 AdderSubtractor_0/fullAdder_2/AND2IN_1/NOT_0/in vdd AdderSubtractor_0/fullAdder_2/AND2IN_1/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1434 AdderSubtractor_0/fullAdder_3/vcin AdderSubtractor_0/fullAdder_2/OR2IN_0/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1435 AdderSubtractor_0/fullAdder_3/vcin AdderSubtractor_0/fullAdder_2/OR2IN_0/NOT_0/in vdd AdderSubtractor_0/fullAdder_2/OR2IN_0/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1436 AdderSubtractor_0/fullAdder_2/OR2IN_0/NOT_0/in AdderSubtractor_0/fullAdder_2/OR2IN_0/vin2 AdderSubtractor_0/fullAdder_2/OR2IN_0/a_0_1# AdderSubtractor_0/fullAdder_2/OR2IN_0/w_n19_n9# CMOSP w=12 l=2
+  ad=72 pd=36 as=48 ps=32
M1437 AdderSubtractor_0/fullAdder_2/OR2IN_0/NOT_0/in AdderSubtractor_0/fullAdder_2/OR2IN_0/vin2 gnd Gnd CMOSN w=4 l=2
+  ad=60 pd=46 as=0 ps=0
M1438 AdderSubtractor_0/fullAdder_2/OR2IN_0/a_0_1# AdderSubtractor_0/fullAdder_2/OR2IN_0/vin1 vdd AdderSubtractor_0/fullAdder_2/OR2IN_0/w_n19_n9# CMOSP w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1439 AdderSubtractor_0/fullAdder_2/OR2IN_0/NOT_0/in AdderSubtractor_0/fullAdder_2/OR2IN_0/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1440 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_0/a_n1_n23# AdderSubtractor_0/fullAdder_3/XOR2IN_1/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1441 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_3/XOR2IN_1/vin1 vdd AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1442 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_3/vcin AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1443 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_3/vcin vdd AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1444 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_1/a_n1_n23# AdderSubtractor_0/fullAdder_3/XOR2IN_1/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1445 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_3/vin1 AdderSubtractor_0/fullAdder_3/XOR2IN_1/vin1 vdd AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1446 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_3/vin1 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_1/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1447 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_3/vin1 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_2/vin2 vdd AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1448 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_2/a_n1_n23# AdderSubtractor_0/fullAdder_3/vcin gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1449 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_3/vin2 AdderSubtractor_0/fullAdder_3/vcin vdd AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1450 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_3/vin2 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_2/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1451 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_3/vin2 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_2/vin2 vdd AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1452 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_3/a_n1_n23# AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_3/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1453 OR2IN_1/vin1 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_3/vin1 vdd AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1454 OR2IN_1/vin1 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_3/vin2 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_3/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1455 OR2IN_1/vin1 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_3/vin2 vdd AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1456 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_0/a_n1_n23# Enable_0/vouta3 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1457 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_2/vin2 Enable_0/vouta3 vdd AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1458 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_2/vin2 AdderSubtractor_0/XOR2IN_3/vout AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1459 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_2/vin2 AdderSubtractor_0/XOR2IN_3/vout vdd AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1460 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_1/a_n1_n23# Enable_0/vouta3 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1461 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_3/vin1 Enable_0/vouta3 vdd AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1462 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_3/vin1 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_1/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1463 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_3/vin1 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_2/vin2 vdd AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1464 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_2/a_n1_n23# AdderSubtractor_0/XOR2IN_3/vout gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1465 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_3/vin2 AdderSubtractor_0/XOR2IN_3/vout vdd AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1466 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_3/vin2 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_2/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1467 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_3/vin2 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_2/vin2 vdd AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1468 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_3/a_n1_n23# AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_3/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1469 AdderSubtractor_0/fullAdder_3/XOR2IN_1/vin1 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_3/vin1 vdd AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1470 AdderSubtractor_0/fullAdder_3/XOR2IN_1/vin1 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_3/vin2 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_3/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1471 AdderSubtractor_0/fullAdder_3/XOR2IN_1/vin1 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_3/vin2 vdd AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1472 AdderSubtractor_0/fullAdder_3/AND2IN_0/NAND2IN_0/a_n1_n23# Enable_0/vouta3 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1473 AdderSubtractor_0/fullAdder_3/AND2IN_0/NOT_0/in Enable_0/vouta3 vdd AdderSubtractor_0/fullAdder_3/AND2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1474 AdderSubtractor_0/fullAdder_3/AND2IN_0/NOT_0/in AdderSubtractor_0/XOR2IN_3/vout AdderSubtractor_0/fullAdder_3/AND2IN_0/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1475 AdderSubtractor_0/fullAdder_3/AND2IN_0/NOT_0/in AdderSubtractor_0/XOR2IN_3/vout vdd AdderSubtractor_0/fullAdder_3/AND2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1476 AdderSubtractor_0/fullAdder_3/OR2IN_0/vin2 AdderSubtractor_0/fullAdder_3/AND2IN_0/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1477 AdderSubtractor_0/fullAdder_3/OR2IN_0/vin2 AdderSubtractor_0/fullAdder_3/AND2IN_0/NOT_0/in vdd AdderSubtractor_0/fullAdder_3/AND2IN_0/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1478 AdderSubtractor_0/fullAdder_3/AND2IN_1/NAND2IN_0/a_n1_n23# AdderSubtractor_0/fullAdder_3/vcin gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1479 AdderSubtractor_0/fullAdder_3/AND2IN_1/NOT_0/in AdderSubtractor_0/fullAdder_3/vcin vdd AdderSubtractor_0/fullAdder_3/AND2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1480 AdderSubtractor_0/fullAdder_3/AND2IN_1/NOT_0/in AdderSubtractor_0/fullAdder_3/XOR2IN_1/vin1 AdderSubtractor_0/fullAdder_3/AND2IN_1/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1481 AdderSubtractor_0/fullAdder_3/AND2IN_1/NOT_0/in AdderSubtractor_0/fullAdder_3/XOR2IN_1/vin1 vdd AdderSubtractor_0/fullAdder_3/AND2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1482 AdderSubtractor_0/fullAdder_3/OR2IN_0/vin1 AdderSubtractor_0/fullAdder_3/AND2IN_1/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1483 AdderSubtractor_0/fullAdder_3/OR2IN_0/vin1 AdderSubtractor_0/fullAdder_3/AND2IN_1/NOT_0/in vdd AdderSubtractor_0/fullAdder_3/AND2IN_1/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1484 vcout AdderSubtractor_0/fullAdder_3/OR2IN_0/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1485 vcout AdderSubtractor_0/fullAdder_3/OR2IN_0/NOT_0/in vdd AdderSubtractor_0/fullAdder_3/OR2IN_0/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1486 AdderSubtractor_0/fullAdder_3/OR2IN_0/NOT_0/in AdderSubtractor_0/fullAdder_3/OR2IN_0/vin2 AdderSubtractor_0/fullAdder_3/OR2IN_0/a_0_1# AdderSubtractor_0/fullAdder_3/OR2IN_0/w_n19_n9# CMOSP w=12 l=2
+  ad=72 pd=36 as=48 ps=32
M1487 AdderSubtractor_0/fullAdder_3/OR2IN_0/NOT_0/in AdderSubtractor_0/fullAdder_3/OR2IN_0/vin2 gnd Gnd CMOSN w=4 l=2
+  ad=60 pd=46 as=0 ps=0
M1488 AdderSubtractor_0/fullAdder_3/OR2IN_0/a_0_1# AdderSubtractor_0/fullAdder_3/OR2IN_0/vin1 vdd AdderSubtractor_0/fullAdder_3/OR2IN_0/w_n19_n9# CMOSP w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1489 AdderSubtractor_0/fullAdder_3/OR2IN_0/NOT_0/in AdderSubtractor_0/fullAdder_3/OR2IN_0/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1490 AdderSubtractor_0/XOR2IN_0/NAND2IN_0/a_n1_n23# Enable_0/voutb0 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1491 AdderSubtractor_0/XOR2IN_0/NAND2IN_2/vin2 Enable_0/voutb0 vdd AdderSubtractor_0/XOR2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1492 AdderSubtractor_0/XOR2IN_0/NAND2IN_2/vin2 OR2IN_0/vin2 AdderSubtractor_0/XOR2IN_0/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1493 AdderSubtractor_0/XOR2IN_0/NAND2IN_2/vin2 OR2IN_0/vin2 vdd AdderSubtractor_0/XOR2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1494 AdderSubtractor_0/XOR2IN_0/NAND2IN_1/a_n1_n23# Enable_0/voutb0 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1495 AdderSubtractor_0/XOR2IN_0/NAND2IN_3/vin1 Enable_0/voutb0 vdd AdderSubtractor_0/XOR2IN_0/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1496 AdderSubtractor_0/XOR2IN_0/NAND2IN_3/vin1 AdderSubtractor_0/XOR2IN_0/NAND2IN_2/vin2 AdderSubtractor_0/XOR2IN_0/NAND2IN_1/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1497 AdderSubtractor_0/XOR2IN_0/NAND2IN_3/vin1 AdderSubtractor_0/XOR2IN_0/NAND2IN_2/vin2 vdd AdderSubtractor_0/XOR2IN_0/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1498 AdderSubtractor_0/XOR2IN_0/NAND2IN_2/a_n1_n23# OR2IN_0/vin2 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1499 AdderSubtractor_0/XOR2IN_0/NAND2IN_3/vin2 OR2IN_0/vin2 vdd AdderSubtractor_0/XOR2IN_0/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1500 AdderSubtractor_0/XOR2IN_0/NAND2IN_3/vin2 AdderSubtractor_0/XOR2IN_0/NAND2IN_2/vin2 AdderSubtractor_0/XOR2IN_0/NAND2IN_2/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1501 AdderSubtractor_0/XOR2IN_0/NAND2IN_3/vin2 AdderSubtractor_0/XOR2IN_0/NAND2IN_2/vin2 vdd AdderSubtractor_0/XOR2IN_0/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1502 AdderSubtractor_0/XOR2IN_0/NAND2IN_3/a_n1_n23# AdderSubtractor_0/XOR2IN_0/NAND2IN_3/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1503 AdderSubtractor_0/XOR2IN_0/vout AdderSubtractor_0/XOR2IN_0/NAND2IN_3/vin1 vdd AdderSubtractor_0/XOR2IN_0/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1504 AdderSubtractor_0/XOR2IN_0/vout AdderSubtractor_0/XOR2IN_0/NAND2IN_3/vin2 AdderSubtractor_0/XOR2IN_0/NAND2IN_3/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1505 AdderSubtractor_0/XOR2IN_0/vout AdderSubtractor_0/XOR2IN_0/NAND2IN_3/vin2 vdd AdderSubtractor_0/XOR2IN_0/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1506 AdderSubtractor_0/XOR2IN_1/NAND2IN_0/a_n1_n23# Enable_0/voutb1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1507 AdderSubtractor_0/XOR2IN_1/NAND2IN_2/vin2 Enable_0/voutb1 vdd AdderSubtractor_0/XOR2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1508 AdderSubtractor_0/XOR2IN_1/NAND2IN_2/vin2 OR2IN_0/vin2 AdderSubtractor_0/XOR2IN_1/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1509 AdderSubtractor_0/XOR2IN_1/NAND2IN_2/vin2 OR2IN_0/vin2 vdd AdderSubtractor_0/XOR2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1510 AdderSubtractor_0/XOR2IN_1/NAND2IN_1/a_n1_n23# Enable_0/voutb1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1511 AdderSubtractor_0/XOR2IN_1/NAND2IN_3/vin1 Enable_0/voutb1 vdd AdderSubtractor_0/XOR2IN_1/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1512 AdderSubtractor_0/XOR2IN_1/NAND2IN_3/vin1 AdderSubtractor_0/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/XOR2IN_1/NAND2IN_1/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1513 AdderSubtractor_0/XOR2IN_1/NAND2IN_3/vin1 AdderSubtractor_0/XOR2IN_1/NAND2IN_2/vin2 vdd AdderSubtractor_0/XOR2IN_1/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1514 AdderSubtractor_0/XOR2IN_1/NAND2IN_2/a_n1_n23# OR2IN_0/vin2 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1515 AdderSubtractor_0/XOR2IN_1/NAND2IN_3/vin2 OR2IN_0/vin2 vdd AdderSubtractor_0/XOR2IN_1/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1516 AdderSubtractor_0/XOR2IN_1/NAND2IN_3/vin2 AdderSubtractor_0/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/XOR2IN_1/NAND2IN_2/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1517 AdderSubtractor_0/XOR2IN_1/NAND2IN_3/vin2 AdderSubtractor_0/XOR2IN_1/NAND2IN_2/vin2 vdd AdderSubtractor_0/XOR2IN_1/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1518 AdderSubtractor_0/XOR2IN_1/NAND2IN_3/a_n1_n23# AdderSubtractor_0/XOR2IN_1/NAND2IN_3/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1519 AdderSubtractor_0/XOR2IN_1/vout AdderSubtractor_0/XOR2IN_1/NAND2IN_3/vin1 vdd AdderSubtractor_0/XOR2IN_1/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1520 AdderSubtractor_0/XOR2IN_1/vout AdderSubtractor_0/XOR2IN_1/NAND2IN_3/vin2 AdderSubtractor_0/XOR2IN_1/NAND2IN_3/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1521 AdderSubtractor_0/XOR2IN_1/vout AdderSubtractor_0/XOR2IN_1/NAND2IN_3/vin2 vdd AdderSubtractor_0/XOR2IN_1/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1522 AdderSubtractor_0/XOR2IN_2/NAND2IN_0/a_n1_n23# Enable_0/voutb2 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1523 AdderSubtractor_0/XOR2IN_2/NAND2IN_2/vin2 Enable_0/voutb2 vdd AdderSubtractor_0/XOR2IN_2/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1524 AdderSubtractor_0/XOR2IN_2/NAND2IN_2/vin2 OR2IN_0/vin2 AdderSubtractor_0/XOR2IN_2/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1525 AdderSubtractor_0/XOR2IN_2/NAND2IN_2/vin2 OR2IN_0/vin2 vdd AdderSubtractor_0/XOR2IN_2/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1526 AdderSubtractor_0/XOR2IN_2/NAND2IN_1/a_n1_n23# Enable_0/voutb2 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1527 AdderSubtractor_0/XOR2IN_2/NAND2IN_3/vin1 Enable_0/voutb2 vdd AdderSubtractor_0/XOR2IN_2/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1528 AdderSubtractor_0/XOR2IN_2/NAND2IN_3/vin1 AdderSubtractor_0/XOR2IN_2/NAND2IN_2/vin2 AdderSubtractor_0/XOR2IN_2/NAND2IN_1/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1529 AdderSubtractor_0/XOR2IN_2/NAND2IN_3/vin1 AdderSubtractor_0/XOR2IN_2/NAND2IN_2/vin2 vdd AdderSubtractor_0/XOR2IN_2/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1530 AdderSubtractor_0/XOR2IN_2/NAND2IN_2/a_n1_n23# OR2IN_0/vin2 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1531 AdderSubtractor_0/XOR2IN_2/NAND2IN_3/vin2 OR2IN_0/vin2 vdd AdderSubtractor_0/XOR2IN_2/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1532 AdderSubtractor_0/XOR2IN_2/NAND2IN_3/vin2 AdderSubtractor_0/XOR2IN_2/NAND2IN_2/vin2 AdderSubtractor_0/XOR2IN_2/NAND2IN_2/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1533 AdderSubtractor_0/XOR2IN_2/NAND2IN_3/vin2 AdderSubtractor_0/XOR2IN_2/NAND2IN_2/vin2 vdd AdderSubtractor_0/XOR2IN_2/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1534 AdderSubtractor_0/XOR2IN_2/NAND2IN_3/a_n1_n23# AdderSubtractor_0/XOR2IN_2/NAND2IN_3/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1535 AdderSubtractor_0/XOR2IN_2/vout AdderSubtractor_0/XOR2IN_2/NAND2IN_3/vin1 vdd AdderSubtractor_0/XOR2IN_2/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1536 AdderSubtractor_0/XOR2IN_2/vout AdderSubtractor_0/XOR2IN_2/NAND2IN_3/vin2 AdderSubtractor_0/XOR2IN_2/NAND2IN_3/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1537 AdderSubtractor_0/XOR2IN_2/vout AdderSubtractor_0/XOR2IN_2/NAND2IN_3/vin2 vdd AdderSubtractor_0/XOR2IN_2/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1538 AdderSubtractor_0/XOR2IN_3/NAND2IN_0/a_n1_n23# Enable_0/voutb3 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1539 AdderSubtractor_0/XOR2IN_3/NAND2IN_2/vin2 Enable_0/voutb3 vdd AdderSubtractor_0/XOR2IN_3/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1540 AdderSubtractor_0/XOR2IN_3/NAND2IN_2/vin2 OR2IN_0/vin2 AdderSubtractor_0/XOR2IN_3/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1541 AdderSubtractor_0/XOR2IN_3/NAND2IN_2/vin2 OR2IN_0/vin2 vdd AdderSubtractor_0/XOR2IN_3/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1542 AdderSubtractor_0/XOR2IN_3/NAND2IN_1/a_n1_n23# Enable_0/voutb3 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1543 AdderSubtractor_0/XOR2IN_3/NAND2IN_3/vin1 Enable_0/voutb3 vdd AdderSubtractor_0/XOR2IN_3/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1544 AdderSubtractor_0/XOR2IN_3/NAND2IN_3/vin1 AdderSubtractor_0/XOR2IN_3/NAND2IN_2/vin2 AdderSubtractor_0/XOR2IN_3/NAND2IN_1/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1545 AdderSubtractor_0/XOR2IN_3/NAND2IN_3/vin1 AdderSubtractor_0/XOR2IN_3/NAND2IN_2/vin2 vdd AdderSubtractor_0/XOR2IN_3/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1546 AdderSubtractor_0/XOR2IN_3/NAND2IN_2/a_n1_n23# OR2IN_0/vin2 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1547 AdderSubtractor_0/XOR2IN_3/NAND2IN_3/vin2 OR2IN_0/vin2 vdd AdderSubtractor_0/XOR2IN_3/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1548 AdderSubtractor_0/XOR2IN_3/NAND2IN_3/vin2 AdderSubtractor_0/XOR2IN_3/NAND2IN_2/vin2 AdderSubtractor_0/XOR2IN_3/NAND2IN_2/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1549 AdderSubtractor_0/XOR2IN_3/NAND2IN_3/vin2 AdderSubtractor_0/XOR2IN_3/NAND2IN_2/vin2 vdd AdderSubtractor_0/XOR2IN_3/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1550 AdderSubtractor_0/XOR2IN_3/NAND2IN_3/a_n1_n23# AdderSubtractor_0/XOR2IN_3/NAND2IN_3/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1551 AdderSubtractor_0/XOR2IN_3/vout AdderSubtractor_0/XOR2IN_3/NAND2IN_3/vin1 vdd AdderSubtractor_0/XOR2IN_3/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1552 AdderSubtractor_0/XOR2IN_3/vout AdderSubtractor_0/XOR2IN_3/NAND2IN_3/vin2 AdderSubtractor_0/XOR2IN_3/NAND2IN_3/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1553 AdderSubtractor_0/XOR2IN_3/vout AdderSubtractor_0/XOR2IN_3/NAND2IN_3/vin2 vdd AdderSubtractor_0/XOR2IN_3/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1554 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_0/a_n1_n23# AdderSubtractor_0/fullAdder_0/XOR2IN_1/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1555 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_0/XOR2IN_1/vin1 vdd AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1556 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_2/vin2 OR2IN_0/vin2 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1557 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_2/vin2 OR2IN_0/vin2 vdd AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1558 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_1/a_n1_n23# AdderSubtractor_0/fullAdder_0/XOR2IN_1/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1559 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_3/vin1 AdderSubtractor_0/fullAdder_0/XOR2IN_1/vin1 vdd AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1560 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_3/vin1 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_1/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1561 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_3/vin1 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_2/vin2 vdd AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1562 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_2/a_n1_n23# OR2IN_0/vin2 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1563 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_3/vin2 OR2IN_0/vin2 vdd AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1564 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_3/vin2 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_2/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1565 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_3/vin2 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_2/vin2 vdd AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1566 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_3/a_n1_n23# AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_3/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1567 OR3IN_0/vin1 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_3/vin1 vdd AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1568 OR3IN_0/vin1 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_3/vin2 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_3/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1569 OR3IN_0/vin1 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_3/vin2 vdd AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1570 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_0/a_n1_n23# Enable_0/vouta0 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1571 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_2/vin2 Enable_0/vouta0 vdd AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1572 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_2/vin2 AdderSubtractor_0/XOR2IN_0/vout AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1573 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_2/vin2 AdderSubtractor_0/XOR2IN_0/vout vdd AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1574 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_1/a_n1_n23# Enable_0/vouta0 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1575 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_3/vin1 Enable_0/vouta0 vdd AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1576 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_3/vin1 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_1/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1577 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_3/vin1 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_2/vin2 vdd AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1578 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_2/a_n1_n23# AdderSubtractor_0/XOR2IN_0/vout gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1579 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_3/vin2 AdderSubtractor_0/XOR2IN_0/vout vdd AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1580 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_3/vin2 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_2/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1581 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_3/vin2 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_2/vin2 vdd AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1582 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_3/a_n1_n23# AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_3/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1583 AdderSubtractor_0/fullAdder_0/XOR2IN_1/vin1 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_3/vin1 vdd AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1584 AdderSubtractor_0/fullAdder_0/XOR2IN_1/vin1 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_3/vin2 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_3/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1585 AdderSubtractor_0/fullAdder_0/XOR2IN_1/vin1 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_3/vin2 vdd AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1586 AdderSubtractor_0/fullAdder_0/AND2IN_0/NAND2IN_0/a_n1_n23# Enable_0/vouta0 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1587 AdderSubtractor_0/fullAdder_0/AND2IN_0/NOT_0/in Enable_0/vouta0 vdd AdderSubtractor_0/fullAdder_0/AND2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1588 AdderSubtractor_0/fullAdder_0/AND2IN_0/NOT_0/in AdderSubtractor_0/XOR2IN_0/vout AdderSubtractor_0/fullAdder_0/AND2IN_0/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1589 AdderSubtractor_0/fullAdder_0/AND2IN_0/NOT_0/in AdderSubtractor_0/XOR2IN_0/vout vdd AdderSubtractor_0/fullAdder_0/AND2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1590 AdderSubtractor_0/fullAdder_0/OR2IN_0/vin2 AdderSubtractor_0/fullAdder_0/AND2IN_0/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1591 AdderSubtractor_0/fullAdder_0/OR2IN_0/vin2 AdderSubtractor_0/fullAdder_0/AND2IN_0/NOT_0/in vdd AdderSubtractor_0/fullAdder_0/AND2IN_0/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1592 AdderSubtractor_0/fullAdder_0/AND2IN_1/NAND2IN_0/a_n1_n23# OR2IN_0/vin2 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1593 AdderSubtractor_0/fullAdder_0/AND2IN_1/NOT_0/in OR2IN_0/vin2 vdd AdderSubtractor_0/fullAdder_0/AND2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1594 AdderSubtractor_0/fullAdder_0/AND2IN_1/NOT_0/in AdderSubtractor_0/fullAdder_0/XOR2IN_1/vin1 AdderSubtractor_0/fullAdder_0/AND2IN_1/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1595 AdderSubtractor_0/fullAdder_0/AND2IN_1/NOT_0/in AdderSubtractor_0/fullAdder_0/XOR2IN_1/vin1 vdd AdderSubtractor_0/fullAdder_0/AND2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1596 AdderSubtractor_0/fullAdder_0/OR2IN_0/vin1 AdderSubtractor_0/fullAdder_0/AND2IN_1/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1597 AdderSubtractor_0/fullAdder_0/OR2IN_0/vin1 AdderSubtractor_0/fullAdder_0/AND2IN_1/NOT_0/in vdd AdderSubtractor_0/fullAdder_0/AND2IN_1/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1598 AdderSubtractor_0/fullAdder_1/vcin AdderSubtractor_0/fullAdder_0/OR2IN_0/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1599 AdderSubtractor_0/fullAdder_1/vcin AdderSubtractor_0/fullAdder_0/OR2IN_0/NOT_0/in vdd AdderSubtractor_0/fullAdder_0/OR2IN_0/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1600 AdderSubtractor_0/fullAdder_0/OR2IN_0/NOT_0/in AdderSubtractor_0/fullAdder_0/OR2IN_0/vin2 AdderSubtractor_0/fullAdder_0/OR2IN_0/a_0_1# AdderSubtractor_0/fullAdder_0/OR2IN_0/w_n19_n9# CMOSP w=12 l=2
+  ad=72 pd=36 as=48 ps=32
M1601 AdderSubtractor_0/fullAdder_0/OR2IN_0/NOT_0/in AdderSubtractor_0/fullAdder_0/OR2IN_0/vin2 gnd Gnd CMOSN w=4 l=2
+  ad=60 pd=46 as=0 ps=0
M1602 AdderSubtractor_0/fullAdder_0/OR2IN_0/a_0_1# AdderSubtractor_0/fullAdder_0/OR2IN_0/vin1 vdd AdderSubtractor_0/fullAdder_0/OR2IN_0/w_n19_n9# CMOSP w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1603 AdderSubtractor_0/fullAdder_0/OR2IN_0/NOT_0/in AdderSubtractor_0/fullAdder_0/OR2IN_0/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1604 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_0/a_n1_n23# AdderSubtractor_0/fullAdder_1/XOR2IN_1/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1605 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_1/XOR2IN_1/vin1 vdd AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1606 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_1/vcin AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1607 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_1/vcin vdd AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1608 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_1/a_n1_n23# AdderSubtractor_0/fullAdder_1/XOR2IN_1/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1609 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_3/vin1 AdderSubtractor_0/fullAdder_1/XOR2IN_1/vin1 vdd AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1610 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_3/vin1 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_1/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1611 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_3/vin1 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_2/vin2 vdd AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1612 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_2/a_n1_n23# AdderSubtractor_0/fullAdder_1/vcin gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1613 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_3/vin2 AdderSubtractor_0/fullAdder_1/vcin vdd AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1614 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_3/vin2 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_2/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1615 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_3/vin2 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_2/vin2 vdd AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1616 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_3/a_n1_n23# AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_3/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1617 OR3IN_1/vin1 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_3/vin1 vdd AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1618 OR3IN_1/vin1 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_3/vin2 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_3/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1619 OR3IN_1/vin1 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_3/vin2 vdd AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1620 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_0/a_n1_n23# Enable_0/vouta1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1621 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_2/vin2 Enable_0/vouta1 vdd AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1622 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_2/vin2 AdderSubtractor_0/XOR2IN_1/vout AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1623 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_2/vin2 AdderSubtractor_0/XOR2IN_1/vout vdd AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1624 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_1/a_n1_n23# Enable_0/vouta1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1625 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_3/vin1 Enable_0/vouta1 vdd AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1626 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_3/vin1 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_1/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1627 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_3/vin1 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_2/vin2 vdd AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1628 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_2/a_n1_n23# AdderSubtractor_0/XOR2IN_1/vout gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1629 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_3/vin2 AdderSubtractor_0/XOR2IN_1/vout vdd AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1630 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_3/vin2 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_2/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1631 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_3/vin2 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_2/vin2 vdd AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1632 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_3/a_n1_n23# AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_3/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1633 AdderSubtractor_0/fullAdder_1/XOR2IN_1/vin1 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_3/vin1 vdd AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1634 AdderSubtractor_0/fullAdder_1/XOR2IN_1/vin1 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_3/vin2 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_3/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1635 AdderSubtractor_0/fullAdder_1/XOR2IN_1/vin1 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_3/vin2 vdd AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1636 AdderSubtractor_0/fullAdder_1/AND2IN_0/NAND2IN_0/a_n1_n23# Enable_0/vouta1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1637 AdderSubtractor_0/fullAdder_1/AND2IN_0/NOT_0/in Enable_0/vouta1 vdd AdderSubtractor_0/fullAdder_1/AND2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1638 AdderSubtractor_0/fullAdder_1/AND2IN_0/NOT_0/in AdderSubtractor_0/XOR2IN_1/vout AdderSubtractor_0/fullAdder_1/AND2IN_0/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1639 AdderSubtractor_0/fullAdder_1/AND2IN_0/NOT_0/in AdderSubtractor_0/XOR2IN_1/vout vdd AdderSubtractor_0/fullAdder_1/AND2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1640 AdderSubtractor_0/fullAdder_1/OR2IN_0/vin2 AdderSubtractor_0/fullAdder_1/AND2IN_0/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1641 AdderSubtractor_0/fullAdder_1/OR2IN_0/vin2 AdderSubtractor_0/fullAdder_1/AND2IN_0/NOT_0/in vdd AdderSubtractor_0/fullAdder_1/AND2IN_0/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1642 AdderSubtractor_0/fullAdder_1/AND2IN_1/NAND2IN_0/a_n1_n23# AdderSubtractor_0/fullAdder_1/vcin gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1643 AdderSubtractor_0/fullAdder_1/AND2IN_1/NOT_0/in AdderSubtractor_0/fullAdder_1/vcin vdd AdderSubtractor_0/fullAdder_1/AND2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1644 AdderSubtractor_0/fullAdder_1/AND2IN_1/NOT_0/in AdderSubtractor_0/fullAdder_1/XOR2IN_1/vin1 AdderSubtractor_0/fullAdder_1/AND2IN_1/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1645 AdderSubtractor_0/fullAdder_1/AND2IN_1/NOT_0/in AdderSubtractor_0/fullAdder_1/XOR2IN_1/vin1 vdd AdderSubtractor_0/fullAdder_1/AND2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1646 AdderSubtractor_0/fullAdder_1/OR2IN_0/vin1 AdderSubtractor_0/fullAdder_1/AND2IN_1/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1647 AdderSubtractor_0/fullAdder_1/OR2IN_0/vin1 AdderSubtractor_0/fullAdder_1/AND2IN_1/NOT_0/in vdd AdderSubtractor_0/fullAdder_1/AND2IN_1/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1648 AdderSubtractor_0/fullAdder_2/vcin AdderSubtractor_0/fullAdder_1/OR2IN_0/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1649 AdderSubtractor_0/fullAdder_2/vcin AdderSubtractor_0/fullAdder_1/OR2IN_0/NOT_0/in vdd AdderSubtractor_0/fullAdder_1/OR2IN_0/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1650 AdderSubtractor_0/fullAdder_1/OR2IN_0/NOT_0/in AdderSubtractor_0/fullAdder_1/OR2IN_0/vin2 AdderSubtractor_0/fullAdder_1/OR2IN_0/a_0_1# AdderSubtractor_0/fullAdder_1/OR2IN_0/w_n19_n9# CMOSP w=12 l=2
+  ad=72 pd=36 as=48 ps=32
M1651 AdderSubtractor_0/fullAdder_1/OR2IN_0/NOT_0/in AdderSubtractor_0/fullAdder_1/OR2IN_0/vin2 gnd Gnd CMOSN w=4 l=2
+  ad=60 pd=46 as=0 ps=0
M1652 AdderSubtractor_0/fullAdder_1/OR2IN_0/a_0_1# AdderSubtractor_0/fullAdder_1/OR2IN_0/vin1 vdd AdderSubtractor_0/fullAdder_1/OR2IN_0/w_n19_n9# CMOSP w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1653 AdderSubtractor_0/fullAdder_1/OR2IN_0/NOT_0/in AdderSubtractor_0/fullAdder_1/OR2IN_0/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
C0 OR2IN_0/vin2 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_2/w_n16_n4# 0.10fF
C1 Comparator_0/NOT_5/out Comparator_0/AND4IN_0/w_n14_n10# 0.15fF
C2 gnd vina2 0.19fF
C3 Decoder_0/AND4Bit_0/AND2IN_0/NOT_0/w_n7_n3# Decoder_0/AND4Bit_0/AND2IN_0/NOT_0/in 0.07fF
C4 AdderSubtractor_0/fullAdder_3/AND2IN_1/NAND2IN_0/w_n16_n4# AdderSubtractor_0/fullAdder_3/AND2IN_1/NOT_0/in 0.08fF
C5 vdd AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_0/w_n16_n4# 0.11fF
C6 gnd Enable_0/voutb2 0.34fF
C7 Enable_1/vouta3 Comparator_0/NOT_2/out 0.06fF
C8 Comparator_0/AND2IN_2/NAND2IN_0/w_n16_n4# Comparator_0/OR4IN_0/vout 0.10fF
C9 Comparator_0/AND2IN_1/NOT_0/w_n7_n3# Comparator_0/AND2IN_1/NOT_0/in 0.07fF
C10 OR3IN_2/w_n19_n9# OR3IN_2/vin3 0.12fF
C11 AdderSubtractor_0/XOR2IN_2/vout AdderSubtractor_0/XOR2IN_2/NAND2IN_3/vin2 0.06fF
C12 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_1/w_n16_n4# AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_2/vin2 0.10fF
C13 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_2/w_n16_n4# AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_2/vin2 0.10fF
C14 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_0/w_n16_n4# vdd 0.11fF
C15 Enable_2/vinEn Enable_2/AND4Bit_0/AND2IN_1/NAND2IN_0/w_n16_n4# 0.10fF
C16 AdderSubtractor_0/XOR2IN_0/NAND2IN_1/w_n16_n4# AdderSubtractor_0/XOR2IN_0/NAND2IN_2/vin2 0.10fF
C17 vina3 Enable_1/AND4Bit_0/AND2IN_3/NAND2IN_0/w_n16_n4# 0.10fF
C18 gnd Enable_1/AND4Bit_0/AND2IN_1/NOT_0/in 0.05fF
C19 Comparator_0/XOR2IN_1/NAND2IN_3/w_n16_n4# Comparator_0/NOT_6/in 0.08fF
C20 Comparator_0/NOT_7/w_n7_n3# Comparator_0/NOT_7/out 0.03fF
C21 Enable_0/voutb3 vdd 0.18fF
C22 vdd Decoder_0/AND4Bit_0/AND2IN_0/NAND2IN_0/w_n16_n4# 0.11fF
C23 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_1/w_n16_n4# AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_2/vin2 0.10fF
C24 AdderSubtractor_0/XOR2IN_3/NAND2IN_3/vin2 vdd 0.08fF
C25 AdderSubtractor_0/XOR2IN_0/NAND2IN_3/w_n16_n4# AdderSubtractor_0/XOR2IN_0/NAND2IN_3/vin1 0.10fF
C26 Enable_2/AND4Bit_1/AND2IN_0/NOT_0/w_n7_n3# vdd 0.06fF
C27 Comparator_0/XOR2IN_2/NAND2IN_3/vin2 Comparator_0/XOR2IN_2/NAND2IN_3/w_n16_n4# 0.10fF
C28 AdderSubtractor_0/fullAdder_3/vcin AdderSubtractor_0/fullAdder_3/XOR2IN_1/vin1 0.26fF
C29 OR3IN_1/NOT_0/in gnd 0.26fF
C30 Enable_1/AND4Bit_0/AND2IN_2/NOT_0/in vdd 0.08fF
C31 Comparator_0/XOR2IN_2/NAND2IN_0/w_n16_n4# Enable_1/voutb2 0.10fF
C32 Enable_1/voutb0 gnd 0.23fF
C33 Comparator_0/XOR2IN_3/NAND2IN_2/w_n16_n4# Comparator_0/XOR2IN_3/NAND2IN_3/vin2 0.08fF
C34 OR2IN_0/vin2 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_0/w_n16_n4# 0.10fF
C35 AdderSubtractor_0/fullAdder_2/OR2IN_0/vin2 AdderSubtractor_0/fullAdder_2/OR2IN_0/vin1 0.11fF
C36 Enable_2/vinEn vdd 0.18fF
C37 Comparator_0/OR4IN_0/NOT_0/w_n7_n3# Comparator_0/OR4IN_0/vout 0.03fF
C38 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_3/vin2 0.06fF
C39 Enable_1/vouta3 Enable_1/voutb3 0.06fF
C40 Comparator_0/XOR2IN_0/NAND2IN_3/vin2 vdd 0.08fF
C41 OR3IN_1/vin2 vcout 0.06fF
C42 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_0/w_n16_n4# AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_2/vin2 0.08fF
C43 AdderSubtractor_0/fullAdder_1/OR2IN_0/NOT_0/w_n7_n3# AdderSubtractor_0/fullAdder_1/OR2IN_0/NOT_0/in 0.07fF
C44 Comparator_0/NOT_7/w_n7_n3# vdd 0.06fF
C45 AdderSubtractor_0/fullAdder_2/OR2IN_0/vin2 AdderSubtractor_0/fullAdder_2/OR2IN_0/w_n19_n9# 0.12fF
C46 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_3/vin2 0.06fF
C47 gnd Enable_0/AND4Bit_0/AND2IN_0/NOT_0/in 0.05fF
C48 Enable_1/AND4Bit_1/AND2IN_1/NOT_0/in vdd 0.08fF
C49 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_3/vin1 0.06fF
C50 Comparator_0/OR4IN_0/vin3 Comparator_0/OR4IN_0/w_n19_n9# 0.12fF
C51 AdderSubtractor_0/fullAdder_2/OR2IN_0/NOT_0/w_n7_n3# AdderSubtractor_0/fullAdder_2/OR2IN_0/NOT_0/in 0.07fF
C52 Comparator_0/AND4IN_1/NOT_0/in Comparator_0/AND4IN_1/w_n14_n10# 0.25fF
C53 AdderSubtractor_0/fullAdder_0/AND2IN_0/NAND2IN_0/w_n16_n4# vdd 0.11fF
C54 AdderSubtractor_0/XOR2IN_3/NAND2IN_3/w_n16_n4# AdderSubtractor_0/XOR2IN_3/NAND2IN_3/vin1 0.10fF
C55 vinb2 Enable_1/AND4Bit_1/AND2IN_2/NAND2IN_0/w_n16_n4# 0.10fF
C56 OR3IN_2/vin2 vcout 0.06fF
C57 Comparator_0/OR4IN_0/vin4 Comparator_0/OR4IN_0/NOT_0/in 0.13fF
C58 Comparator_0/NOT_5/out Enable_1/vouta2 0.06fF
C59 Comparator_0/XOR2IN_1/NAND2IN_3/vin1 gnd 0.13fF
C60 Comparator_0/NOT_6/out Comparator_0/AND4IN_0/NOT_0/in 0.06fF
C61 OR3IN_2/NOT_0/in OR3IN_2/w_n19_n9# 0.05fF
C62 OR3IN_0/vin2 OR3IN_0/vin1 0.14fF
C63 Enable_1/voutb2 gnd 0.29fF
C64 gnd AdderSubtractor_0/fullAdder_1/XOR2IN_1/vin1 0.52fF
C65 gnd AdderSubtractor_0/fullAdder_3/OR2IN_0/NOT_0/in 0.11fF
C66 AdderSubtractor_0/fullAdder_3/AND2IN_0/NOT_0/in AdderSubtractor_0/fullAdder_3/AND2IN_0/NOT_0/w_n7_n3# 0.07fF
C67 AdderSubtractor_0/fullAdder_1/vcin AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_2/w_n16_n4# 0.10fF
C68 vdd AdderSubtractor_0/fullAdder_0/AND2IN_1/NOT_0/w_n7_n3# 0.06fF
C69 OR2IN_0/vout vinb0 0.06fF
C70 AND4Bit_0/AND2IN_3/NAND2IN_0/w_n16_n4# Enable_2/voutb3 0.10fF
C71 Comparator_0/NOT_4/out Comparator_0/NOT_4/w_n7_n3# 0.03fF
C72 vout0 OR3IN_0/NOT_0/w_n7_n3# 0.03fF
C73 Enable_0/vouta2 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_0/w_n16_n4# 0.10fF
C74 Enable_0/AND4Bit_0/AND2IN_1/NAND2IN_0/w_n16_n4# Enable_0/AND4Bit_0/AND2IN_1/NOT_0/in 0.08fF
C75 gnd OR2IN_1/vin1 0.12fF
C76 AdderSubtractor_0/XOR2IN_0/vout AdderSubtractor_0/fullAdder_0/AND2IN_0/NAND2IN_0/w_n16_n4# 0.10fF
C77 Enable_0/voutb2 AdderSubtractor_0/XOR2IN_2/NAND2IN_1/w_n16_n4# 0.10fF
C78 AND4Bit_0/AND2IN_0/NOT_0/in gnd 0.05fF
C79 Enable_0/AND4Bit_0/AND2IN_1/NOT_0/in gnd 0.05fF
C80 Comparator_0/XOR2IN_0/NAND2IN_3/w_n16_n4# Comparator_0/XOR2IN_0/NAND2IN_3/vin1 0.10fF
C81 Comparator_0/AND5IN_0/NOT_0/in Comparator_0/NOT_3/out 0.06fF
C82 AdderSubtractor_0/fullAdder_0/AND2IN_1/NOT_0/w_n7_n3# AdderSubtractor_0/fullAdder_0/OR2IN_0/vin1 0.03fF
C83 gnd Enable_1/AND4Bit_1/AND2IN_0/NOT_0/in 0.05fF
C84 Enable_1/vouta1 Enable_1/AND4Bit_0/AND2IN_1/NOT_0/w_n7_n3# 0.03fF
C85 gnd Comparator_0/NOT_4/out 0.45fF
C86 vout0 gnd 0.07fF
C87 Enable_0/vouta3 OR2IN_0/vin2 0.13fF
C88 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_0/w_n16_n4# AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_2/vin2 0.08fF
C89 Enable_2/AND4Bit_0/AND2IN_2/NAND2IN_0/w_n16_n4# Enable_2/AND4Bit_0/AND2IN_2/NOT_0/in 0.08fF
C90 vinb0 vinb3 0.19fF
C91 Comparator_0/AND5IN_0/NOT_0/in Comparator_0/AND5IN_0/w_n26_1# 0.24fF
C92 OR3IN_1/w_n19_n9# OR3IN_1/vin1 0.16fF
C93 vina3 vinb2 0.19fF
C94 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_0/w_n16_n4# AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_2/vin2 0.08fF
C95 Enable_0/AND4Bit_1/AND2IN_0/NOT_0/w_n7_n3# vdd 0.06fF
C96 Enable_1/voutb0 Comparator_0/XOR2IN_0/NAND2IN_2/vin2 0.39fF
C97 AdderSubtractor_0/fullAdder_3/OR2IN_0/vin2 AdderSubtractor_0/fullAdder_3/AND2IN_0/NOT_0/w_n7_n3# 0.03fF
C98 Enable_0/AND4Bit_0/AND2IN_3/NAND2IN_0/w_n16_n4# vdd 0.11fF
C99 Comparator_0/XOR2IN_1/NAND2IN_3/vin2 Comparator_0/NOT_6/in 0.06fF
C100 AdderSubtractor_0/fullAdder_3/XOR2IN_1/vin1 vdd 0.21fF
C101 Enable_1/vouta3 gnd 0.53fF
C102 OR2IN_0/vin2 AdderSubtractor_0/XOR2IN_3/NAND2IN_2/w_n16_n4# 0.10fF
C103 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_1/w_n16_n4# AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_3/vin1 0.08fF
C104 OR3IN_1/NOT_0/in OR3IN_1/NOT_0/w_n7_n3# 0.07fF
C105 AdderSubtractor_0/fullAdder_3/OR2IN_0/vin2 AdderSubtractor_0/fullAdder_3/OR2IN_0/NOT_0/in 0.08fF
C106 Enable_2/AND4Bit_0/AND2IN_2/NOT_0/w_n7_n3# vdd 0.06fF
C107 Comparator_0/NOT_0/out vdd 0.06fF
C108 OR3IN_1/vin3 vcout 0.06fF
C109 Comparator_0/NOT_2/out vdd 0.06fF
C110 Comparator_0/XOR2IN_3/NAND2IN_3/w_n16_n4# Comparator_0/XOR2IN_3/NAND2IN_3/vin1 0.10fF
C111 AdderSubtractor_0/XOR2IN_3/NAND2IN_1/w_n16_n4# AdderSubtractor_0/XOR2IN_3/NAND2IN_3/vin1 0.08fF
C112 Decoder_0/NOT_1/w_n7_n3# vdd 0.06fF
C113 Enable_0/AND4Bit_0/AND2IN_3/NAND2IN_0/w_n16_n4# Enable_0/AND4Bit_0/AND2IN_3/NOT_0/in 0.08fF
C114 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_2/w_n16_n4# vdd 0.11fF
C115 AND4Bit_0/AND2IN_3/NOT_0/w_n7_n3# vdd 0.06fF
C116 Comparator_0/XOR2IN_2/NAND2IN_3/vin1 vdd 0.43fF
C117 gnd AdderSubtractor_0/fullAdder_3/vcin 0.48fF
C118 Enable_2/AND4Bit_1/AND2IN_1/NOT_0/w_n7_n3# vdd 0.06fF
C119 Enable_1/vinEn vinb1 0.13fF
C120 Comparator_0/AND2IN_1/NAND2IN_0/w_n16_n4# Enable_1/vinEn 0.10fF
C121 Comparator_0/AND2IN_0/NOT_0/in vdd 0.08fF
C122 gnd AdderSubtractor_0/fullAdder_1/AND2IN_1/NOT_0/in 0.05fF
C123 Decoder_0/AND4Bit_0/AND2IN_2/NOT_0/w_n7_n3# vdd 0.06fF
C124 Enable_1/vinEn Enable_1/AND4Bit_1/AND2IN_3/NOT_0/in 0.06fF
C125 Enable_1/voutb3 vdd 0.18fF
C126 gnd Enable_0/vouta3 0.53fF
C127 Enable_1/voutb1 Comparator_0/XOR2IN_1/NAND2IN_2/vin2 0.39fF
C128 AdderSubtractor_0/fullAdder_0/XOR2IN_1/vin1 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_3/w_n16_n4# 0.08fF
C129 gnd AdderSubtractor_0/fullAdder_2/AND2IN_1/NOT_0/in 0.05fF
C130 OR2IN_0/vin2 AdderSubtractor_0/XOR2IN_2/NAND2IN_2/vin2 0.39fF
C131 AdderSubtractor_0/XOR2IN_0/NAND2IN_3/vin2 AdderSubtractor_0/XOR2IN_0/NAND2IN_3/w_n16_n4# 0.10fF
C132 AdderSubtractor_0/fullAdder_2/vcin AdderSubtractor_0/fullAdder_1/OR2IN_0/NOT_0/w_n7_n3# 0.03fF
C133 OR3IN_0/NOT_0/w_n7_n3# OR3IN_0/NOT_0/in 0.07fF
C134 AdderSubtractor_0/XOR2IN_0/vout AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_2/w_n16_n4# 0.10fF
C135 Decoder_0/NOT_0/w_n7_n3# Decoder_0/NOT_0/out 0.03fF
C136 gnd Enable_2/AND4Bit_0/AND2IN_3/NOT_0/in 0.05fF
C137 Enable_2/AND4Bit_0/AND2IN_2/NOT_0/w_n7_n3# Enable_2/vouta2 0.03fF
C138 OR2IN_0/vin2 vdd 0.32fF
C139 Enable_2/vinEn Enable_2/AND4Bit_1/AND2IN_1/NAND2IN_0/w_n16_n4# 0.10fF
C140 Comparator_0/AND2IN_1/NOT_0/in Comparator_0/AND4IN_0/vout 0.06fF
C141 Comparator_0/NOT_0/out Comparator_0/AND2IN_0/NAND2IN_0/w_n16_n4# 0.10fF
C142 Enable_1/AND4Bit_0/AND2IN_2/NAND2IN_0/w_n16_n4# Enable_1/AND4Bit_0/AND2IN_2/NOT_0/in 0.08fF
C143 Comparator_0/AND3IN_0/NOT_0/w_n7_n3# Comparator_0/AND3IN_0/NOT_0/in 0.07fF
C144 Enable_2/AND4Bit_1/AND2IN_0/NOT_0/in Enable_2/AND4Bit_1/AND2IN_0/NAND2IN_0/w_n16_n4# 0.08fF
C145 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_2/vin2 vdd 0.08fF
C146 AdderSubtractor_0/XOR2IN_0/NAND2IN_2/vin2 vdd 0.08fF
C147 Comparator_0/XOR2IN_2/NAND2IN_0/w_n16_n4# vdd 0.11fF
C148 gnd OR3IN_0/NOT_0/in 0.26fF
C149 AdderSubtractor_0/fullAdder_3/AND2IN_1/NOT_0/in vdd 0.08fF
C150 Enable_2/AND4Bit_0/AND2IN_3/NAND2IN_0/w_n16_n4# Enable_2/AND4Bit_0/AND2IN_3/NOT_0/in 0.08fF
C151 AdderSubtractor_0/fullAdder_3/vcin AdderSubtractor_0/fullAdder_3/OR2IN_0/vin2 0.06fF
C152 OR3IN_2/vin3 AND4Bit_0/AND2IN_2/NOT_0/w_n7_n3# 0.03fF
C153 OR3IN_0/w_n19_n9# OR3IN_0/vin3 0.12fF
C154 Enable_1/vinEn Enable_1/AND4Bit_0/AND2IN_3/NAND2IN_0/w_n16_n4# 0.10fF
C155 Enable_0/voutb3 AdderSubtractor_0/XOR2IN_3/NAND2IN_0/w_n16_n4# 0.10fF
C156 AdderSubtractor_0/fullAdder_3/XOR2IN_1/vin1 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_3/w_n16_n4# 0.08fF
C157 Comparator_0/XOR2IN_3/NAND2IN_1/w_n16_n4# Comparator_0/XOR2IN_3/NAND2IN_3/vin1 0.08fF
C158 gnd Enable_2/AND4Bit_1/AND2IN_2/NOT_0/in 0.05fF
C159 OR2IN_1/vin2 OR2IN_1/vin1 0.11fF
C160 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_3/vin1 0.06fF
C161 Comparator_0/AND2IN_0/NAND2IN_0/w_n16_n4# Comparator_0/AND2IN_0/NOT_0/in 0.08fF
C162 vdd AdderSubtractor_0/fullAdder_0/OR2IN_0/NOT_0/w_n7_n3# 0.06fF
C163 Enable_0/AND4Bit_0/AND2IN_2/NOT_0/w_n7_n3# vdd 0.06fF
C164 Comparator_0/NOT_7/out gnd 0.20fF
C165 Enable_2/AND4Bit_1/AND2IN_3/NOT_0/in vdd 0.08fF
C166 Comparator_0/NOT_5/w_n7_n3# Comparator_0/NOT_5/out 0.03fF
C167 gnd AdderSubtractor_0/fullAdder_1/AND2IN_0/NOT_0/in 0.05fF
C168 Enable_1/vinEn Enable_1/AND4Bit_1/AND2IN_2/NAND2IN_0/w_n16_n4# 0.10fF
C169 Enable_1/vouta1 Comparator_0/XOR2IN_1/NAND2IN_1/w_n16_n4# 0.10fF
C170 gnd AdderSubtractor_0/fullAdder_2/AND2IN_0/NOT_0/in 0.05fF
C171 vinb3 Enable_2/AND4Bit_1/AND2IN_3/NAND2IN_0/w_n16_n4# 0.10fF
C172 Comparator_0/NOT_4/w_n7_n3# vdd 0.06fF
C173 gnd AdderSubtractor_0/XOR2IN_2/NAND2IN_2/vin2 0.19fF
C174 Enable_2/AND4Bit_1/AND2IN_1/NOT_0/w_n7_n3# Enable_2/voutb1 0.03fF
C175 OR3IN_0/NOT_0/w_n7_n3# vdd 0.06fF
C176 Comparator_0/NOT_5/out Enable_1/vouta0 0.19fF
C177 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_3/vcin 0.39fF
C178 Comparator_0/AND2IN_3/NAND2IN_0/w_n16_n4# vdd 0.11fF
C179 AdderSubtractor_0/XOR2IN_1/NAND2IN_3/w_n16_n4# AdderSubtractor_0/XOR2IN_1/vout 0.08fF
C180 Enable_0/AND4Bit_0/AND2IN_1/NAND2IN_0/w_n16_n4# vdd 0.11fF
C181 Enable_0/AND4Bit_0/AND2IN_0/NOT_0/w_n7_n3# Enable_0/AND4Bit_0/AND2IN_0/NOT_0/in 0.07fF
C182 vina1 OR2IN_0/vout 0.06fF
C183 Enable_0/AND4Bit_1/AND2IN_1/NOT_0/w_n7_n3# vdd 0.06fF
C184 Enable_2/AND4Bit_1/AND2IN_2/NAND2IN_0/w_n16_n4# Enable_2/AND4Bit_1/AND2IN_2/NOT_0/in 0.08fF
C185 gnd vdd 3.53fF
C186 Decoder_0/AND4Bit_0/AND2IN_3/NAND2IN_0/w_n16_n4# Decoder_0/AND4Bit_0/AND2IN_3/NOT_0/in 0.08fF
C187 AdderSubtractor_0/XOR2IN_3/NAND2IN_2/w_n16_n4# AdderSubtractor_0/XOR2IN_3/NAND2IN_2/vin2 0.10fF
C188 Enable_1/vinEn Comparator_0/AND2IN_3/NOT_0/in 0.06fF
C189 gnd AdderSubtractor_0/fullAdder_1/OR2IN_0/vin2 0.27fF
C190 Decoder_0/AND4Bit_0/AND2IN_0/NAND2IN_0/w_n16_n4# Decoder_0/NOT_1/out 0.10fF
C191 Enable_0/vouta2 OR2IN_0/vin2 0.13fF
C192 gnd AdderSubtractor_0/fullAdder_0/OR2IN_0/vin1 0.26fF
C193 AdderSubtractor_0/XOR2IN_2/NAND2IN_3/w_n16_n4# vdd 0.11fF
C194 AdderSubtractor_0/fullAdder_3/AND2IN_0/NOT_0/in vdd 0.08fF
C195 Enable_2/AND4Bit_0/AND2IN_3/NAND2IN_0/w_n16_n4# vdd 0.11fF
C196 Comparator_0/NOT_5/in Comparator_0/NOT_4/out 0.07fF
C197 vina1 vinb3 0.19fF
C198 gnd AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_3/vin1 0.06fF
C199 AdderSubtractor_0/fullAdder_0/XOR2IN_1/vin1 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_3/vin2 0.06fF
C200 Comparator_0/NOT_1/out Comparator_0/NOT_2/out 5.84fF
C201 OR3IN_2/vin3 OR3IN_2/vin2 0.14fF
C202 Comparator_0/OR4IN_0/vin2 Comparator_0/OR4IN_0/w_n19_n9# 0.12fF
C203 Enable_1/vinEn vina3 0.13fF
C204 gnd Enable_0/AND4Bit_0/AND2IN_3/NOT_0/in 0.05fF
C205 Comparator_0/OR4IN_0/vin2 Comparator_0/OR4IN_0/vin3 0.18fF
C206 gnd AdderSubtractor_0/XOR2IN_1/NAND2IN_3/vin2 0.06fF
C207 gnd AdderSubtractor_0/XOR2IN_0/vout 0.28fF
C208 Enable_1/AND4Bit_1/AND2IN_0/NOT_0/in Enable_1/AND4Bit_1/AND2IN_0/NAND2IN_0/w_n16_n4# 0.08fF
C209 Enable_2/AND4Bit_1/AND2IN_2/NAND2IN_0/w_n16_n4# vdd 0.11fF
C210 Comparator_0/XOR2IN_1/NAND2IN_2/w_n16_n4# vdd 0.11fF
C211 Comparator_0/XOR2IN_0/NAND2IN_2/w_n16_n4# Comparator_0/XOR2IN_0/NAND2IN_2/vin2 0.10fF
C212 AdderSubtractor_0/XOR2IN_1/vout AdderSubtractor_0/fullAdder_1/AND2IN_0/NOT_0/in 0.06fF
C213 Enable_1/AND4Bit_0/AND2IN_3/NAND2IN_0/w_n16_n4# Enable_1/AND4Bit_0/AND2IN_3/NOT_0/in 0.08fF
C214 Comparator_0/NOT_5/out Comparator_0/AND4IN_1/w_n14_n10# 0.15fF
C215 vinSel0 Decoder_0/NOT_1/out 0.50fF
C216 vdd AdderSubtractor_0/fullAdder_1/OR2IN_0/vin1 0.06fF
C217 Enable_1/vinEn Enable_1/AND4Bit_0/AND2IN_0/NOT_0/in 0.06fF
C218 Enable_0/AND4Bit_0/AND2IN_2/NOT_0/w_n7_n3# Enable_0/vouta2 0.03fF
C219 gnd AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_2/vin2 0.19fF
C220 AdderSubtractor_0/fullAdder_3/OR2IN_0/vin2 vdd 0.06fF
C221 vout2 OR3IN_2/NOT_0/w_n7_n3# 0.03fF
C222 AdderSubtractor_0/fullAdder_2/OR2IN_0/vin1 vdd 0.06fF
C223 AdderSubtractor_0/fullAdder_2/vcin AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_2/vin2 0.39fF
C224 vdd AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_3/vin1 0.43fF
C225 AdderSubtractor_0/XOR2IN_2/vout AdderSubtractor_0/fullAdder_2/AND2IN_0/NOT_0/in 0.06fF
C226 Enable_1/vinEn vinb2 0.13fF
C227 gnd Enable_0/AND4Bit_1/AND2IN_2/NOT_0/in 0.05fF
C228 Enable_1/voutb3 Comparator_0/NOT_1/out 0.06fF
C229 OR2IN_0/vout Enable_0/AND4Bit_1/AND2IN_3/NAND2IN_0/w_n16_n4# 0.10fF
C230 AdderSubtractor_0/fullAdder_1/OR2IN_0/vin2 AdderSubtractor_0/fullAdder_1/OR2IN_0/vin1 0.11fF
C231 vdd AdderSubtractor_0/fullAdder_1/OR2IN_0/w_n19_n9# 0.09fF
C232 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_3/vin1 vdd 0.43fF
C233 gnd Enable_2/vouta2 0.14fF
C234 Comparator_0/NOT_5/out Comparator_0/NOT_3/out 0.19fF
C235 OR3IN_1/w_n19_n9# OR3IN_1/vin2 0.12fF
C236 Enable_0/vouta1 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_0/w_n16_n4# 0.10fF
C237 OR2IN_0/vin2 AdderSubtractor_0/fullAdder_0/OR2IN_0/vin2 0.06fF
C238 AdderSubtractor_0/fullAdder_3/XOR2IN_1/vin1 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_3/vin2 0.06fF
C239 Enable_1/vouta0 Enable_1/AND4Bit_0/AND2IN_0/NOT_0/w_n7_n3# 0.03fF
C240 Comparator_0/NOT_4/in Comparator_0/NOT_4/w_n7_n3# 0.07fF
C241 AdderSubtractor_0/fullAdder_2/OR2IN_0/w_n19_n9# vdd 0.09fF
C242 Enable_0/AND4Bit_1/AND2IN_3/NOT_0/in vdd 0.08fF
C243 vdd AdderSubtractor_0/XOR2IN_1/vout 0.20fF
C244 AdderSubtractor_0/XOR2IN_3/NAND2IN_2/vin2 vdd 0.08fF
C245 Comparator_0/NOT_5/out Comparator_0/AND5IN_0/w_n26_1# 0.12fF
C246 AdderSubtractor_0/fullAdder_1/OR2IN_0/vin2 AdderSubtractor_0/fullAdder_1/OR2IN_0/w_n19_n9# 0.12fF
C247 AdderSubtractor_0/XOR2IN_2/NAND2IN_1/w_n16_n4# AdderSubtractor_0/XOR2IN_2/NAND2IN_2/vin2 0.10fF
C248 Enable_2/vouta3 vdd 0.15fF
C249 AdderSubtractor_0/XOR2IN_2/vout vdd 0.20fF
C250 Enable_0/AND4Bit_1/AND2IN_3/NAND2IN_0/w_n16_n4# vinb3 0.10fF
C251 gnd Enable_0/vouta2 0.53fF
C252 Enable_1/voutb0 Enable_1/vouta3 19.55fF
C253 Comparator_0/NOT_4/in gnd 0.07fF
C254 Comparator_0/XOR2IN_3/NAND2IN_2/w_n16_n4# Comparator_0/XOR2IN_3/NAND2IN_2/vin2 0.10fF
C255 vdd Decoder_0/AND4Bit_0/AND2IN_1/NOT_0/in 0.08fF
C256 gnd Enable_2/voutb1 0.14fF
C257 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_1/w_n16_n4# AdderSubtractor_0/fullAdder_3/XOR2IN_1/vin1 0.10fF
C258 Comparator_0/OR4IN_0/NOT_0/w_n7_n3# Comparator_0/OR4IN_0/NOT_0/in 0.07fF
C259 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_2/w_n16_n4# AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_3/vin2 0.08fF
C260 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_2/vin2 vdd 0.08fF
C261 AdderSubtractor_0/XOR2IN_2/NAND2IN_1/w_n16_n4# vdd 0.11fF
C262 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_3/vin2 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_3/w_n16_n4# 0.10fF
C263 Comparator_0/XOR2IN_0/NAND2IN_2/vin2 vdd 0.08fF
C264 Enable_1/AND4Bit_1/AND2IN_2/NAND2IN_0/w_n16_n4# Enable_1/AND4Bit_1/AND2IN_2/NOT_0/in 0.08fF
C265 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_3/w_n16_n4# AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_3/vin1 0.10fF
C266 OR3IN_2/NOT_0/in OR3IN_2/vin2 0.08fF
C267 Enable_2/voutb2 vdd 0.19fF
C268 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_2/w_n16_n4# AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_3/vin2 0.08fF
C269 OR3IN_2/vin3 OR3IN_1/vin3 0.06fF
C270 AdderSubtractor_0/XOR2IN_1/NAND2IN_3/vin2 AdderSubtractor_0/XOR2IN_1/vout 0.06fF
C271 Enable_1/vouta2 Comparator_0/NOT_0/out 0.06fF
C272 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_3/vin1 0.06fF
C273 AdderSubtractor_0/XOR2IN_2/NAND2IN_2/vin2 AdderSubtractor_0/XOR2IN_2/NAND2IN_3/vin2 0.06fF
C274 OR3IN_1/NOT_0/w_n7_n3# vdd 0.06fF
C275 Enable_0/voutb2 Enable_0/vouta3 0.06fF
C276 Enable_1/vouta2 Comparator_0/NOT_2/out 0.06fF
C277 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_3/vin1 vdd 0.43fF
C278 Enable_2/AND4Bit_0/AND2IN_0/NOT_0/in vdd 0.08fF
C279 Enable_0/voutb1 OR2IN_0/vin2 0.06fF
C280 Comparator_0/AND2IN_2/NOT_0/in Comparator_0/OR4IN_0/vout 0.06fF
C281 vout3 vdd 0.08fF
C282 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_1/w_n16_n4# AdderSubtractor_0/fullAdder_0/XOR2IN_1/vin1 0.10fF
C283 AdderSubtractor_0/XOR2IN_2/NAND2IN_3/vin2 vdd 0.08fF
C284 gnd AdderSubtractor_0/fullAdder_0/OR2IN_0/vin2 0.27fF
C285 OR2IN_1/vin2 vdd 0.06fF
C286 vinb1 vinb0 2.82fF
C287 OR2IN_0/vin2 AdderSubtractor_0/XOR2IN_3/NAND2IN_0/w_n16_n4# 0.10fF
C288 Enable_0/AND4Bit_1/AND2IN_2/NAND2IN_0/w_n16_n4# vdd 0.11fF
C289 Enable_0/AND4Bit_1/AND2IN_0/NOT_0/in Enable_0/AND4Bit_1/AND2IN_0/NAND2IN_0/w_n16_n4# 0.08fF
C290 Enable_1/vouta2 Enable_1/voutb3 0.06fF
C291 Enable_1/voutb2 Enable_1/vouta3 0.06fF
C292 Comparator_0/AND2IN_1/NAND2IN_0/w_n16_n4# Comparator_0/AND2IN_1/NOT_0/in 0.08fF
C293 Comparator_0/NOR2IN_0/w_n19_n9# OR3IN_0/vin2 0.16fF
C294 vdd AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_3/vin2 0.08fF
C295 AND4Bit_0/AND2IN_3/NOT_0/in Enable_2/voutb3 0.06fF
C296 Comparator_0/AND5IN_0/NOT_0/in Comparator_0/NOT_6/out 0.06fF
C297 OR3IN_2/vin2 Comparator_0/NOR2IN_0/vout 0.41fF
C298 Enable_2/vinEn Enable_2/AND4Bit_0/AND2IN_2/NOT_0/in 0.06fF
C299 OR2IN_0/NOT_0/in OR2IN_0/vin2 0.08fF
C300 Decoder_0/NOT_1/w_n7_n3# Decoder_0/NOT_1/out 0.03fF
C301 Decoder_0/AND4Bit_0/AND2IN_2/NOT_0/in vdd 0.08fF
C302 AdderSubtractor_0/fullAdder_3/vcin AdderSubtractor_0/fullAdder_3/AND2IN_1/NAND2IN_0/w_n16_n4# 0.10fF
C303 Comparator_0/NOT_1/out gnd 2.09fF
C304 gnd AdderSubtractor_0/XOR2IN_3/NAND2IN_3/vin1 0.13fF
C305 AdderSubtractor_0/fullAdder_0/AND2IN_1/NOT_0/w_n7_n3# AdderSubtractor_0/fullAdder_0/AND2IN_1/NOT_0/in 0.07fF
C306 vinb3 Enable_2/vinEn 0.20fF
C307 Comparator_0/XOR2IN_2/NAND2IN_1/w_n16_n4# Comparator_0/XOR2IN_2/NAND2IN_2/vin2 0.10fF
C308 Enable_0/vouta2 AdderSubtractor_0/XOR2IN_2/vout 0.27fF
C309 Enable_2/vouta3 Enable_2/voutb1 0.06fF
C310 AND4Bit_0/AND2IN_0/NAND2IN_0/w_n16_n4# Enable_2/voutb0 0.10fF
C311 Comparator_0/NOT_3/out Comparator_0/NOT_3/w_n7_n3# 0.03fF
C312 OR3IN_1/w_n19_n9# OR3IN_1/vin3 0.12fF
C313 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_0/w_n16_n4# vdd 0.11fF
C314 Enable_1/vouta3 Comparator_0/NOT_4/out 0.06fF
C315 Comparator_0/OR4IN_0/vin4 gnd 0.19fF
C316 Enable_2/vinEn Enable_2/AND4Bit_1/AND2IN_1/NOT_0/in 0.06fF
C317 Comparator_0/XOR2IN_0/NAND2IN_3/vin1 gnd 0.13fF
C318 AdderSubtractor_0/fullAdder_2/OR2IN_0/vin2 vdd 0.06fF
C319 Comparator_0/NOT_5/out Enable_1/vouta1 0.13fF
C320 Enable_1/voutb0 Comparator_0/XOR2IN_0/NAND2IN_2/w_n16_n4# 0.10fF
C321 AdderSubtractor_0/XOR2IN_3/vout AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_2/vin2 0.39fF
C322 Comparator_0/NOT_5/in vdd 0.15fF
C323 Enable_1/vouta2 Comparator_0/XOR2IN_2/NAND2IN_0/w_n16_n4# 0.10fF
C324 Enable_1/AND4Bit_1/AND2IN_3/NOT_0/w_n7_n3# vdd 0.06fF
C325 Enable_0/AND4Bit_1/AND2IN_1/NOT_0/w_n7_n3# Enable_0/voutb1 0.03fF
C326 AdderSubtractor_0/fullAdder_1/XOR2IN_1/vin1 AdderSubtractor_0/fullAdder_1/AND2IN_1/NOT_0/in 0.06fF
C327 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_3/w_n16_n4# OR3IN_0/vin1 0.08fF
C328 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_3/vin2 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_3/w_n16_n4# 0.10fF
C329 gnd Enable_0/voutb1 0.34fF
C330 Comparator_0/XOR2IN_2/NAND2IN_2/vin2 Comparator_0/XOR2IN_2/NAND2IN_3/vin2 0.06fF
C331 Enable_1/voutb1 gnd 0.29fF
C332 OR2IN_1/NOT_0/in OR2IN_1/w_n19_n9# 0.05fF
C333 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_3/vin2 0.06fF
C334 AdderSubtractor_0/fullAdder_0/AND2IN_0/NOT_0/in AdderSubtractor_0/fullAdder_0/AND2IN_0/NAND2IN_0/w_n16_n4# 0.08fF
C335 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_3/vin2 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_3/w_n16_n4# 0.10fF
C336 Enable_0/AND4Bit_1/AND2IN_2/NAND2IN_0/w_n16_n4# Enable_0/AND4Bit_1/AND2IN_2/NOT_0/in 0.08fF
C337 Enable_0/voutb2 vdd 0.35fF
C338 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_3/w_n16_n4# AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_3/vin1 0.10fF
C339 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_0/w_n16_n4# AdderSubtractor_0/XOR2IN_0/vout 0.10fF
C340 Enable_1/AND4Bit_1/AND2IN_0/NAND2IN_0/w_n16_n4# vdd 0.11fF
C341 Decoder_0/AND4Bit_0/AND2IN_3/NOT_0/in vinSel1 0.06fF
C342 Decoder_0/AND4Bit_0/AND2IN_3/NAND2IN_0/w_n16_n4# vinSel0 0.10fF
C343 Enable_1/voutb2 Comparator_0/NOT_1/w_n7_n3# 0.07fF
C344 Enable_1/AND4Bit_0/AND2IN_1/NOT_0/in vdd 0.08fF
C345 Enable_0/AND4Bit_0/AND2IN_0/NOT_0/w_n7_n3# vdd 0.06fF
C346 Comparator_0/NOT_6/w_n7_n3# vdd 0.06fF
C347 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_3/w_n16_n4# AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_3/vin1 0.10fF
C348 OR2IN_0/NOT_0/in gnd 0.11fF
C349 Enable_1/voutb0 vdd 0.25fF
C350 AdderSubtractor_0/XOR2IN_3/NAND2IN_2/vin2 AdderSubtractor_0/XOR2IN_3/NAND2IN_3/vin1 0.06fF
C351 OR2IN_0/vout Enable_0/AND4Bit_0/AND2IN_3/NAND2IN_0/w_n16_n4# 0.10fF
C352 OR3IN_0/w_n19_n9# OR3IN_0/vin1 0.16fF
C353 AdderSubtractor_0/fullAdder_3/OR2IN_0/NOT_0/w_n7_n3# vcout 0.03fF
C354 Enable_1/voutb1 Comparator_0/XOR2IN_1/NAND2IN_2/w_n16_n4# 0.10fF
C355 OR2IN_0/vin2 AdderSubtractor_0/XOR2IN_2/NAND2IN_2/w_n16_n4# 0.10fF
C356 vinb1 Enable_1/AND4Bit_1/AND2IN_1/NAND2IN_0/w_n16_n4# 0.10fF
C357 Enable_1/vouta2 gnd 0.53fF
C358 gnd AdderSubtractor_0/fullAdder_1/OR2IN_0/NOT_0/in 0.11fF
C359 OR3IN_0/vin2 vcout 0.06fF
C360 Enable_0/vouta0 AdderSubtractor_0/fullAdder_0/AND2IN_0/NAND2IN_0/w_n16_n4# 0.10fF
C361 gnd AdderSubtractor_0/fullAdder_2/OR2IN_0/NOT_0/in 0.11fF
C362 Enable_0/AND4Bit_0/AND2IN_0/NOT_0/in vdd 0.08fF
C363 AND4Bit_0/AND2IN_3/NAND2IN_0/w_n16_n4# Enable_2/vouta3 0.10fF
C364 gnd OR3IN_1/vin1 0.12fF
C365 AdderSubtractor_0/fullAdder_3/AND2IN_1/NAND2IN_0/w_n16_n4# vdd 0.14fF
C366 Enable_2/AND4Bit_0/AND2IN_2/NOT_0/w_n7_n3# Enable_2/AND4Bit_0/AND2IN_2/NOT_0/in 0.07fF
C367 gnd OR3IN_2/vin1 0.12fF
C368 Enable_0/AND4Bit_0/AND2IN_2/NAND2IN_0/w_n16_n4# vina2 0.10fF
C369 Enable_2/AND4Bit_1/AND2IN_0/NOT_0/w_n7_n3# Enable_2/voutb0 0.03fF
C370 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_2/w_n16_n4# vdd 0.11fF
C371 gnd Decoder_0/NOT_1/out 0.28fF
C372 OR2IN_0/vin2 Enable_0/vouta1 0.13fF
C373 AdderSubtractor_0/XOR2IN_0/NAND2IN_1/w_n16_n4# vdd 0.11fF
C374 Comparator_0/XOR2IN_1/NAND2IN_3/vin1 vdd 0.43fF
C375 Comparator_0/XOR2IN_0/NAND2IN_2/vin2 Comparator_0/XOR2IN_0/NAND2IN_3/vin1 0.06fF
C376 vina3 vinb0 1.48fF
C377 AdderSubtractor_0/fullAdder_3/AND2IN_0/NOT_0/w_n7_n3# vdd 0.09fF
C378 AdderSubtractor_0/fullAdder_3/vcin Enable_0/vouta3 0.06fF
C379 OR2IN_0/vin2 AdderSubtractor_0/XOR2IN_0/NAND2IN_0/w_n16_n4# 0.10fF
C380 Comparator_0/AND3IN_0/NOT_0/in Comparator_0/AND3IN_0/w_n14_n10# 0.19fF
C381 vinb0 Enable_2/AND4Bit_1/AND2IN_0/NAND2IN_0/w_n16_n4# 0.10fF
C382 AdderSubtractor_0/XOR2IN_3/NAND2IN_0/w_n16_n4# AdderSubtractor_0/XOR2IN_3/NAND2IN_2/vin2 0.08fF
C383 vina0 Enable_1/AND4Bit_0/AND2IN_0/NAND2IN_0/w_n16_n4# 0.10fF
C384 Comparator_0/AND2IN_3/NOT_0/w_n7_n3# vdd 0.06fF
C385 gnd AND4Bit_0/AND2IN_2/NOT_0/in 0.05fF
C386 Enable_1/voutb2 vdd 0.25fF
C387 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_1/w_n16_n4# AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_3/vin1 0.08fF
C388 vdd AdderSubtractor_0/fullAdder_1/XOR2IN_1/vin1 0.21fF
C389 AdderSubtractor_0/fullAdder_1/vcin AdderSubtractor_0/fullAdder_0/OR2IN_0/NOT_0/w_n7_n3# 0.03fF
C390 OR2IN_0/vin2 AdderSubtractor_0/XOR2IN_1/NAND2IN_2/vin2 0.39fF
C391 AdderSubtractor_0/XOR2IN_0/NAND2IN_2/vin2 AdderSubtractor_0/XOR2IN_0/NAND2IN_0/w_n16_n4# 0.08fF
C392 Enable_1/vouta0 Comparator_0/NOT_0/out 0.06fF
C393 OR2IN_1/vin1 vdd 0.08fF
C394 Comparator_0/AND3IN_0/w_n14_n10# Comparator_0/NOT_5/out 0.15fF
C395 Enable_1/vouta0 Comparator_0/NOT_2/out 0.06fF
C396 Comparator_0/AND4IN_0/NOT_0/w_n7_n3# vdd 0.06fF
C397 vinb0 vinb2 0.19fF
C398 AND4Bit_0/AND2IN_0/NOT_0/in vdd 0.08fF
C399 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_0/w_n16_n4# vdd 0.11fF
C400 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_1/w_n16_n4# AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_3/vin1 0.08fF
C401 Enable_0/AND4Bit_0/AND2IN_1/NOT_0/in vdd 0.08fF
C402 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_3/vin2 OR3IN_0/vin1 0.06fF
C403 Comparator_0/AND2IN_2/NOT_0/w_n7_n3# vdd 0.06fF
C404 Enable_1/AND4Bit_1/AND2IN_0/NOT_0/in vdd 0.08fF
C405 OR2IN_0/vout OR2IN_0/vin2 0.06fF
C406 Enable_2/AND4Bit_1/AND2IN_1/NOT_0/w_n7_n3# Enable_2/AND4Bit_1/AND2IN_1/NOT_0/in 0.07fF
C407 Comparator_0/NOT_4/out vdd 0.12fF
C408 vout0 vdd 0.24fF
C409 AdderSubtractor_0/fullAdder_1/OR2IN_0/NOT_0/in AdderSubtractor_0/fullAdder_1/OR2IN_0/w_n19_n9# 0.05fF
C410 Comparator_0/XOR2IN_3/NAND2IN_2/vin2 Comparator_0/XOR2IN_3/NAND2IN_3/vin1 0.06fF
C411 vina1 vinb1 0.19fF
C412 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_2/w_n16_n4# vdd 0.11fF
C413 AND4Bit_0/AND2IN_0/NOT_0/in AND4Bit_0/AND2IN_0/NOT_0/w_n7_n3# 0.07fF
C414 AdderSubtractor_0/fullAdder_2/OR2IN_0/NOT_0/in AdderSubtractor_0/fullAdder_2/OR2IN_0/w_n19_n9# 0.05fF
C415 Comparator_0/AND2IN_0/NOT_0/w_n7_n3# Comparator_0/OR4IN_0/vin1 0.03fF
C416 Comparator_0/XOR2IN_1/NAND2IN_0/w_n16_n4# vdd 0.11fF
C417 gnd AdderSubtractor_0/fullAdder_1/vcin 0.48fF
C418 Enable_2/AND4Bit_0/AND2IN_1/NOT_0/w_n7_n3# vdd 0.06fF
C419 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_1/w_n16_n4# 0.10fF
C420 Enable_1/vouta0 Enable_1/voutb3 0.06fF
C421 Enable_1/vouta3 vdd 0.28fF
C422 gnd Enable_0/vouta1 0.53fF
C423 gnd AdderSubtractor_0/fullAdder_0/AND2IN_1/NOT_0/in 0.05fF
C424 Enable_1/vinEn Enable_1/AND4Bit_0/AND2IN_3/NOT_0/in 0.06fF
C425 Decoder_0/NOT_0/out Decoder_0/AND4Bit_0/AND2IN_1/NAND2IN_0/w_n16_n4# 0.10fF
C426 Enable_1/AND4Bit_0/AND2IN_2/NOT_0/w_n7_n3# Enable_1/AND4Bit_0/AND2IN_2/NOT_0/in 0.07fF
C427 gnd AdderSubtractor_0/XOR2IN_1/NAND2IN_2/vin2 0.19fF
C428 Comparator_0/NOT_2/out Comparator_0/AND4IN_1/w_n14_n10# 0.15fF
C429 Comparator_0/NOT_0/out Comparator_0/NOT_0/w_n7_n3# 0.03fF
C430 Enable_1/vinEn Enable_1/AND4Bit_1/AND2IN_2/NOT_0/in 0.06fF
C431 Comparator_0/XOR2IN_3/NAND2IN_0/w_n16_n4# Comparator_0/XOR2IN_3/NAND2IN_2/vin2 0.08fF
C432 AdderSubtractor_0/fullAdder_3/vcin vdd 0.12fF
C433 OR2IN_0/NOT_0/w_n7_n3# vdd 0.06fF
C434 Enable_0/AND4Bit_0/AND2IN_1/NAND2IN_0/w_n16_n4# OR2IN_0/vout 0.10fF
C435 vina0 OR2IN_0/vout 0.06fF
C436 vdd AdderSubtractor_0/fullAdder_1/AND2IN_1/NOT_0/in 0.08fF
C437 Comparator_0/NOT_2/out Comparator_0/NOT_3/out 9.15fF
C438 Comparator_0/NOT_5/out Comparator_0/AND4IN_0/NOT_0/in 0.06fF
C439 gnd OR2IN_0/vout 0.65fF
C440 Enable_0/vouta3 vdd 0.28fF
C441 AdderSubtractor_0/fullAdder_2/AND2IN_1/NOT_0/in vdd 0.08fF
C442 vina2 Enable_1/AND4Bit_0/AND2IN_2/NAND2IN_0/w_n16_n4# 0.10fF
C443 Enable_0/AND4Bit_1/AND2IN_0/NAND2IN_0/w_n16_n4# vinb0 0.10fF
C444 Enable_1/vinEn Enable_1/AND4Bit_0/AND2IN_1/NAND2IN_0/w_n16_n4# 0.10fF
C445 Comparator_0/OR4IN_0/vin1 Comparator_0/OR4IN_0/w_n19_n9# 0.16fF
C446 gnd Enable_2/AND4Bit_0/AND2IN_2/NOT_0/in 0.05fF
C447 AND4Bit_0/AND2IN_2/NOT_0/in Enable_2/voutb2 0.06fF
C448 Enable_0/voutb1 Enable_0/voutb2 4.04fF
C449 AdderSubtractor_0/XOR2IN_1/NAND2IN_3/w_n16_n4# vdd 0.11fF
C450 OR2IN_0/vin2 Enable_0/vouta0 0.06fF
C451 vina0 vinb3 0.19fF
C452 gnd AdderSubtractor_0/fullAdder_2/vcin 0.48fF
C453 AND4Bit_0/AND2IN_3/NOT_0/w_n7_n3# AND4Bit_0/AND2IN_3/NOT_0/in 0.07fF
C454 Comparator_0/NOT_4/in Comparator_0/NOT_4/out 0.06fF
C455 Enable_2/AND4Bit_0/AND2IN_0/NOT_0/w_n7_n3# Enable_2/AND4Bit_0/AND2IN_0/NOT_0/in 0.07fF
C456 Enable_1/vouta3 Comparator_0/AND2IN_0/NAND2IN_0/w_n16_n4# 0.10fF
C457 AdderSubtractor_0/fullAdder_1/vcin AdderSubtractor_0/XOR2IN_1/vout 0.06fF
C458 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_3/vin2 OR3IN_1/vin1 0.06fF
C459 gnd vinb3 0.19fF
C460 Enable_1/voutb3 Comparator_0/NOT_0/w_n7_n3# 0.07fF
C461 Comparator_0/NOT_1/w_n7_n3# vdd 0.06fF
C462 AdderSubtractor_0/XOR2IN_3/NAND2IN_2/w_n16_n4# vdd 0.11fF
C463 Enable_2/AND4Bit_0/AND2IN_3/NOT_0/in vdd 0.08fF
C464 AdderSubtractor_0/XOR2IN_3/vout AdderSubtractor_0/fullAdder_3/AND2IN_0/NAND2IN_0/w_n16_n4# 0.10fF
C465 OR2IN_0/w_n19_n9# OR2IN_0/vin1 0.16fF
C466 OR3IN_0/vin3 gnd 0.19fF
C467 Enable_0/vouta1 AdderSubtractor_0/XOR2IN_1/vout 0.27fF
C468 gnd AdderSubtractor_0/fullAdder_0/AND2IN_0/NOT_0/in 0.05fF
C469 Enable_1/AND4Bit_1/AND2IN_1/NOT_0/w_n7_n3# Enable_1/AND4Bit_1/AND2IN_1/NOT_0/in 0.07fF
C470 vinSel1 vinSel0 0.13fF
C471 AdderSubtractor_0/fullAdder_3/AND2IN_1/NOT_0/w_n7_n3# AdderSubtractor_0/fullAdder_3/OR2IN_0/vin1 0.03fF
C472 Enable_1/voutb3 Comparator_0/NOT_3/out 0.06fF
C473 AdderSubtractor_0/fullAdder_2/OR2IN_0/vin2 AdderSubtractor_0/fullAdder_2/AND2IN_0/NOT_0/w_n7_n3# 0.03fF
C474 gnd Enable_2/AND4Bit_1/AND2IN_1/NOT_0/in 0.05fF
C475 Enable_1/voutb0 Enable_1/voutb1 16.28fF
C476 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_2/w_n16_n4# AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_2/vin2 0.10fF
C477 Comparator_0/XOR2IN_0/NAND2IN_2/w_n16_n4# vdd 0.11fF
C478 Enable_1/vouta0 gnd 0.53fF
C479 AdderSubtractor_0/XOR2IN_1/NAND2IN_3/vin2 AdderSubtractor_0/XOR2IN_1/NAND2IN_3/w_n16_n4# 0.10fF
C480 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_1/w_n16_n4# AdderSubtractor_0/fullAdder_2/XOR2IN_1/vin1 0.10fF
C481 AdderSubtractor_0/fullAdder_2/OR2IN_0/vin2 AdderSubtractor_0/fullAdder_2/OR2IN_0/NOT_0/in 0.08fF
C482 Enable_2/AND4Bit_1/AND2IN_2/NOT_0/in vdd 0.08fF
C483 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_2/w_n16_n4# AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_2/vin2 0.10fF
C484 Comparator_0/OR4IN_0/NOT_0/in Comparator_0/OR4IN_0/w_n19_n9# 0.05fF
C485 Comparator_0/OR4IN_0/vin3 Comparator_0/OR4IN_0/NOT_0/in 0.09fF
C486 AdderSubtractor_0/XOR2IN_2/NAND2IN_2/w_n16_n4# AdderSubtractor_0/XOR2IN_2/NAND2IN_3/vin2 0.08fF
C487 Comparator_0/NOT_7/out vdd 0.06fF
C488 vdd AdderSubtractor_0/fullAdder_1/AND2IN_0/NOT_0/in 0.08fF
C489 vina1 vina3 0.19fF
C490 Enable_2/AND4Bit_0/AND2IN_1/NAND2IN_0/w_n16_n4# vdd 0.11fF
C491 OR2IN_0/vout Enable_0/AND4Bit_1/AND2IN_3/NOT_0/in 0.06fF
C492 Comparator_0/AND5IN_0/NOT_0/w_n7_n3# vdd 0.06fF
C493 AdderSubtractor_0/fullAdder_2/AND2IN_0/NOT_0/in vdd 0.08fF
C494 AdderSubtractor_0/XOR2IN_2/NAND2IN_2/vin2 vdd 0.08fF
C495 Enable_1/voutb2 Enable_1/AND4Bit_1/AND2IN_2/NOT_0/w_n7_n3# 0.03fF
C496 Enable_0/AND4Bit_0/AND2IN_2/NOT_0/w_n7_n3# Enable_0/AND4Bit_0/AND2IN_2/NOT_0/in 0.07fF
C497 vinb1 Enable_2/vinEn 0.19fF
C498 Comparator_0/NOT_1/out Comparator_0/NOT_4/out 0.06fF
C499 Enable_2/AND4Bit_1/AND2IN_3/NOT_0/w_n7_n3# Enable_2/voutb3 0.03fF
C500 gnd Enable_0/vouta0 0.53fF
C501 Comparator_0/NOT_6/in gnd 0.07fF
C502 Enable_0/AND4Bit_1/AND2IN_0/NOT_0/w_n7_n3# Enable_0/voutb0 0.03fF
C503 Enable_1/voutb0 Enable_1/vouta2 0.06fF
C504 vina1 vinb2 0.19fF
C505 AdderSubtractor_0/fullAdder_2/vcin AdderSubtractor_0/XOR2IN_2/vout 0.06fF
C506 Comparator_0/AND4IN_0/w_n14_n10# Comparator_0/NOT_4/out 0.15fF
C507 AdderSubtractor_0/XOR2IN_1/NAND2IN_1/w_n16_n4# vdd 0.11fF
C508 Enable_1/vouta3 Enable_1/AND4Bit_0/AND2IN_3/NOT_0/w_n7_n3# 0.03fF
C509 Enable_1/voutb1 Enable_1/voutb2 13.11fF
C510 Comparator_0/XOR2IN_3/NAND2IN_3/vin2 gnd 0.06fF
C511 OR3IN_1/vin2 gnd 0.19fF
C512 vdd AdderSubtractor_0/fullAdder_1/OR2IN_0/vin2 0.06fF
C513 Enable_1/vinEn vinb0 0.13fF
C514 Enable_1/vouta1 Comparator_0/NOT_0/out 0.06fF
C515 Enable_1/vouta3 Comparator_0/NOT_1/out 0.06fF
C516 vdd AdderSubtractor_0/fullAdder_0/OR2IN_0/vin1 0.06fF
C517 gnd Enable_0/AND4Bit_0/AND2IN_2/NOT_0/in 0.05fF
C518 Comparator_0/AND4IN_0/vout gnd 0.14fF
C519 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_3/vin1 vdd 0.43fF
C520 AND4Bit_0/AND2IN_0/NOT_0/w_n7_n3# vdd 0.06fF
C521 Enable_1/AND4Bit_0/AND2IN_0/NOT_0/w_n7_n3# Enable_1/AND4Bit_0/AND2IN_0/NOT_0/in 0.07fF
C522 Comparator_0/XOR2IN_0/NAND2IN_3/w_n16_n4# Comparator_0/NOT_7/in 0.08fF
C523 OR3IN_0/w_n19_n9# OR3IN_0/vin2 0.12fF
C524 OR3IN_2/vin2 gnd 0.26fF
C525 AdderSubtractor_0/fullAdder_1/XOR2IN_1/vin1 AdderSubtractor_0/fullAdder_1/AND2IN_1/NAND2IN_0/w_n16_n4# 0.10fF
C526 vdd AdderSubtractor_0/fullAdder_0/OR2IN_0/w_n19_n9# 0.09fF
C527 gnd AND4Bit_0/AND2IN_3/NOT_0/in 0.05fF
C528 AdderSubtractor_0/XOR2IN_3/vout AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_2/w_n16_n4# 0.10fF
C529 Enable_0/AND4Bit_0/AND2IN_3/NOT_0/in vdd 0.08fF
C530 AdderSubtractor_0/XOR2IN_1/NAND2IN_3/vin2 vdd 0.08fF
C531 Comparator_0/NOT_3/out gnd 0.20fF
C532 Comparator_0/XOR2IN_1/NAND2IN_3/vin2 Comparator_0/XOR2IN_1/NAND2IN_3/w_n16_n4# 0.10fF
C533 AdderSubtractor_0/XOR2IN_0/vout vdd 0.20fF
C534 Enable_0/AND4Bit_1/AND2IN_1/NOT_0/w_n7_n3# Enable_0/AND4Bit_1/AND2IN_1/NOT_0/in 0.07fF
C535 gnd Enable_2/voutb0 0.14fF
C536 Comparator_0/XOR2IN_1/NAND2IN_0/w_n16_n4# Enable_1/voutb1 0.10fF
C537 AdderSubtractor_0/fullAdder_0/OR2IN_0/vin1 AdderSubtractor_0/fullAdder_0/OR2IN_0/w_n19_n9# 0.16fF
C538 gnd Enable_0/AND4Bit_1/AND2IN_1/NOT_0/in 0.05fF
C539 Comparator_0/XOR2IN_2/NAND2IN_2/w_n16_n4# Comparator_0/XOR2IN_2/NAND2IN_3/vin2 0.08fF
C540 OR2IN_0/vin2 AdderSubtractor_0/XOR2IN_2/NAND2IN_0/w_n16_n4# 0.10fF
C541 OR2IN_0/vout Enable_0/AND4Bit_1/AND2IN_2/NAND2IN_0/w_n16_n4# 0.10fF
C542 gnd Enable_2/vouta1 0.14fF
C543 Enable_1/vouta2 Enable_1/voutb2 0.06fF
C544 Enable_1/voutb1 Enable_1/vouta3 0.10fF
C545 Enable_1/vouta1 Enable_1/voutb3 0.06fF
C546 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_2/vin2 vdd 0.08fF
C547 vina0 Enable_0/AND4Bit_0/AND2IN_0/NAND2IN_0/w_n16_n4# 0.10fF
C548 Enable_0/AND4Bit_1/AND2IN_2/NOT_0/in vdd 0.08fF
C549 gnd AdderSubtractor_0/XOR2IN_2/NAND2IN_3/vin1 0.13fF
C550 OR2IN_1/w_n19_n9# OR2IN_1/vin2 0.12fF
C551 gnd AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_2/vin2 0.19fF
C552 Enable_2/vouta2 vdd 0.19fF
C553 Enable_0/AND4Bit_0/AND2IN_2/NAND2IN_0/w_n16_n4# vdd 0.11fF
C554 Comparator_0/AND2IN_0/NAND2IN_0/w_n16_n4# vdd 0.11fF
C555 Comparator_0/XOR2IN_3/NAND2IN_3/w_n16_n4# Comparator_0/NOT_5/in 0.08fF
C556 Enable_0/voutb0 OR2IN_0/vin2 0.06fF
C557 Enable_1/vouta2 Comparator_0/NOT_4/out 0.06fF
C558 AdderSubtractor_0/XOR2IN_2/NAND2IN_3/w_n16_n4# AdderSubtractor_0/XOR2IN_2/NAND2IN_3/vin1 0.10fF
C559 Comparator_0/NOT_1/w_n7_n3# Comparator_0/NOT_1/out 0.03fF
C560 OR3IN_2/vin1 OR2IN_1/vin1 7.39fF
C561 Enable_0/vouta2 vdd 0.32fF
C562 Enable_0/vouta3 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_1/w_n16_n4# 0.10fF
C563 Comparator_0/NOT_4/in vdd 0.15fF
C564 Enable_2/voutb1 vdd 0.19fF
C565 Enable_0/voutb1 Enable_0/vouta3 0.06fF
C566 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_3/w_n16_n4# vdd 0.11fF
C567 Enable_1/vouta2 Enable_1/vouta3 25.14fF
C568 AdderSubtractor_0/fullAdder_2/vcin AdderSubtractor_0/fullAdder_2/OR2IN_0/vin2 0.06fF
C569 vina2 OR2IN_0/vout 0.06fF
C570 gnd OR3IN_1/vin3 0.27fF
C571 Enable_1/vinEn Enable_1/AND4Bit_1/AND2IN_1/NAND2IN_0/w_n16_n4# 0.10fF
C572 OR2IN_0/vin2 AdderSubtractor_0/fullAdder_0/AND2IN_1/NAND2IN_0/w_n16_n4# 0.10fF
C573 OR2IN_0/NOT_0/in OR2IN_0/NOT_0/w_n7_n3# 0.07fF
C574 Enable_2/vouta3 Enable_2/voutb0 0.06fF
C575 AdderSubtractor_0/fullAdder_1/AND2IN_1/NAND2IN_0/w_n16_n4# AdderSubtractor_0/fullAdder_1/AND2IN_1/NOT_0/in 0.08fF
C576 vina3 Enable_2/vinEn 0.19fF
C577 Comparator_0/NOT_5/w_n7_n3# Comparator_0/NOT_5/in 0.07fF
C578 vina2 vinb3 0.19fF
C579 Enable_2/vinEn Enable_2/AND4Bit_1/AND2IN_0/NAND2IN_0/w_n16_n4# 0.10fF
C580 AdderSubtractor_0/fullAdder_2/AND2IN_1/NAND2IN_0/w_n16_n4# AdderSubtractor_0/fullAdder_2/AND2IN_1/NOT_0/in 0.08fF
C581 Comparator_0/NOT_7/out Comparator_0/AND4IN_0/w_n14_n10# 0.15fF
C582 AdderSubtractor_0/fullAdder_0/OR2IN_0/vin2 vdd 0.06fF
C583 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_1/w_n16_n4# AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_2/vin2 0.10fF
C584 Enable_2/vinEn Enable_2/AND4Bit_0/AND2IN_1/NOT_0/in 0.06fF
C585 AdderSubtractor_0/fullAdder_1/vcin AdderSubtractor_0/fullAdder_1/XOR2IN_1/vin1 0.26fF
C586 Comparator_0/XOR2IN_0/NAND2IN_3/vin2 Comparator_0/NOT_7/in 0.06fF
C587 gnd Enable_0/voutb0 0.34fF
C588 AND4Bit_0/AND2IN_0/NAND2IN_0/w_n16_n4# Enable_2/vouta0 0.10fF
C589 OR2IN_0/vin2 AdderSubtractor_0/XOR2IN_1/NAND2IN_2/w_n16_n4# 0.10fF
C590 vinb2 Enable_2/vinEn 0.19fF
C591 Enable_1/AND4Bit_0/AND2IN_3/NOT_0/w_n7_n3# vdd 0.06fF
C592 Comparator_0/AND4IN_1/NOT_0/w_n7_n3# vdd 0.06fF
C593 Enable_1/vouta1 gnd 0.53fF
C594 Comparator_0/NOT_7/w_n7_n3# Comparator_0/NOT_7/in 0.07fF
C595 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_3/vin2 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_2/w_n16_n4# 0.08fF
C596 AdderSubtractor_0/fullAdder_0/OR2IN_0/vin2 AdderSubtractor_0/fullAdder_0/OR2IN_0/vin1 0.11fF
C597 Enable_2/vouta2 Enable_2/voutb1 0.06fF
C598 Comparator_0/NOT_1/out vdd 0.06fF
C599 Comparator_0/AND5IN_0/NOT_0/w_n7_n3# Comparator_0/OR4IN_0/vin4 0.03fF
C600 AdderSubtractor_0/XOR2IN_3/NAND2IN_3/vin1 vdd 0.43fF
C601 Enable_0/AND4Bit_0/AND2IN_0/NOT_0/in OR2IN_0/vout 0.06fF
C602 Comparator_0/XOR2IN_2/NAND2IN_3/w_n16_n4# Comparator_0/XOR2IN_2/NAND2IN_3/vin1 0.10fF
C603 gnd vinSel1 0.20fF
C604 Enable_0/vouta0 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_0/w_n16_n4# 0.10fF
C605 AdderSubtractor_0/XOR2IN_2/NAND2IN_1/w_n16_n4# AdderSubtractor_0/XOR2IN_2/NAND2IN_3/vin1 0.08fF
C606 Comparator_0/OR4IN_0/vin2 Comparator_0/OR4IN_0/vin1 0.14fF
C607 AdderSubtractor_0/fullAdder_0/OR2IN_0/vin2 AdderSubtractor_0/fullAdder_0/OR2IN_0/w_n19_n9# 0.12fF
C608 Comparator_0/AND4IN_0/w_n14_n10# vdd 0.25fF
C609 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_3/vin2 0.06fF
C610 AdderSubtractor_0/fullAdder_3/XOR2IN_1/vin1 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_0/w_n16_n4# 0.10fF
C611 Enable_1/AND4Bit_1/AND2IN_2/NOT_0/w_n7_n3# vdd 0.06fF
C612 Enable_2/AND4Bit_1/AND2IN_1/NAND2IN_0/w_n16_n4# vdd 0.11fF
C613 AND4Bit_0/AND2IN_3/NAND2IN_0/w_n16_n4# vdd 0.11fF
C614 Comparator_0/OR4IN_0/vin4 vdd 0.12fF
C615 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_3/vin1 0.06fF
C616 AdderSubtractor_0/fullAdder_0/OR2IN_0/NOT_0/w_n7_n3# AdderSubtractor_0/fullAdder_0/OR2IN_0/NOT_0/in 0.07fF
C617 Comparator_0/XOR2IN_0/NAND2IN_3/vin1 vdd 0.43fF
C618 Comparator_0/AND2IN_0/NOT_0/w_n7_n3# Comparator_0/AND2IN_0/NOT_0/in 0.07fF
C619 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_1/w_n16_n4# vdd 0.11fF
C620 Enable_1/voutb0 Enable_1/vouta0 0.06fF
C621 Enable_1/AND4Bit_0/AND2IN_2/NAND2IN_0/w_n16_n4# vdd 0.11fF
C622 Comparator_0/XOR2IN_3/NAND2IN_3/vin2 Comparator_0/NOT_5/in 0.06fF
C623 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_3/vin1 0.06fF
C624 OR3IN_2/vin3 vcout 0.06fF
C625 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_0/w_n16_n4# vdd 0.11fF
C626 vina1 Enable_1/vinEn 0.13fF
C627 Enable_0/voutb1 vdd 0.35fF
C628 Enable_1/voutb1 vdd 0.25fF
C629 Enable_0/voutb1 AdderSubtractor_0/XOR2IN_1/NAND2IN_1/w_n16_n4# 0.10fF
C630 Enable_0/AND4Bit_1/AND2IN_3/NOT_0/w_n7_n3# Enable_0/voutb3 0.03fF
C631 AdderSubtractor_0/fullAdder_1/AND2IN_0/NOT_0/in AdderSubtractor_0/fullAdder_1/AND2IN_0/NOT_0/w_n7_n3# 0.07fF
C632 Enable_0/AND4Bit_0/AND2IN_0/NOT_0/w_n7_n3# Enable_0/vouta0 0.03fF
C633 Comparator_0/NOR2IN_0/w_n19_n9# Comparator_0/NOR2IN_0/vout 0.05fF
C634 OR3IN_2/w_n19_n9# vdd 0.10fF
C635 Enable_0/AND4Bit_0/AND2IN_1/NOT_0/in OR2IN_0/vout 0.06fF
C636 Comparator_0/NOT_6/w_n7_n3# Comparator_0/NOT_6/in 0.07fF
C637 gnd AdderSubtractor_0/fullAdder_0/OR2IN_0/NOT_0/in 0.11fF
C638 AdderSubtractor_0/XOR2IN_3/NAND2IN_0/w_n16_n4# vdd 0.11fF
C639 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_3/vin2 vdd 0.08fF
C640 Comparator_0/OR4IN_0/vin2 Comparator_0/OR4IN_0/NOT_0/in 0.08fF
C641 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_3/vin2 0.06fF
C642 Enable_0/AND4Bit_0/AND2IN_3/NAND2IN_0/w_n16_n4# vina3 0.10fF
C643 vdd AdderSubtractor_0/fullAdder_1/AND2IN_1/NAND2IN_0/w_n16_n4# 0.14fF
C644 AdderSubtractor_0/fullAdder_2/AND2IN_0/NOT_0/in AdderSubtractor_0/fullAdder_2/AND2IN_0/NOT_0/w_n7_n3# 0.07fF
C645 Enable_2/AND4Bit_1/AND2IN_0/NOT_0/w_n7_n3# Enable_2/AND4Bit_1/AND2IN_0/NOT_0/in 0.07fF
C646 OR2IN_1/w_n19_n9# OR2IN_1/vin1 0.16fF
C647 gnd OR3IN_0/vin1 0.12fF
C648 Comparator_0/NOT_0/out Comparator_0/NOT_6/out 0.06fF
C649 vina0 vinb1 0.19fF
C650 AdderSubtractor_0/fullAdder_2/AND2IN_1/NAND2IN_0/w_n16_n4# vdd 0.14fF
C651 Comparator_0/NOT_6/out Comparator_0/NOT_2/out 0.06fF
C652 vout3 OR3IN_1/vin3 0.06fF
C653 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_0/w_n16_n4# AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_2/vin2 0.08fF
C654 gnd vinb1 0.19fF
C655 Enable_2/vinEn Enable_2/AND4Bit_1/AND2IN_0/NOT_0/in 0.06fF
C656 Comparator_0/NOT_5/out Comparator_0/AND4IN_1/NOT_0/in 0.06fF
C657 OR3IN_1/NOT_0/in OR3IN_1/vin2 0.08fF
C658 Decoder_0/AND4Bit_0/AND2IN_0/NOT_0/in Decoder_0/NOT_0/out 0.06fF
C659 OR3IN_0/vin3 OR2IN_1/vin1 0.07fF
C660 vdd AdderSubtractor_0/fullAdder_1/AND2IN_0/NOT_0/w_n7_n3# 0.09fF
C661 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_1/w_n16_n4# vdd 0.11fF
C662 gnd Enable_1/AND4Bit_1/AND2IN_3/NOT_0/in 0.05fF
C663 AND4Bit_0/AND2IN_1/NAND2IN_0/w_n16_n4# vdd 0.11fF
C664 Enable_1/voutb3 Comparator_0/XOR2IN_3/NAND2IN_2/vin2 0.39fF
C665 Enable_1/vouta0 Enable_1/voutb2 0.06fF
C666 AdderSubtractor_0/fullAdder_2/AND2IN_0/NOT_0/w_n7_n3# vdd 0.09fF
C667 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_0/w_n16_n4# AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_2/vin2 0.08fF
C668 Enable_1/vouta2 vdd 0.32fF
C669 Comparator_0/XOR2IN_2/NAND2IN_1/w_n16_n4# Comparator_0/XOR2IN_2/NAND2IN_3/vin1 0.08fF
C670 AdderSubtractor_0/fullAdder_1/OR2IN_0/vin2 AdderSubtractor_0/fullAdder_1/AND2IN_0/NOT_0/w_n7_n3# 0.03fF
C671 AdderSubtractor_0/fullAdder_2/vcin AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_2/w_n16_n4# 0.10fF
C672 Enable_1/voutb0 Enable_1/AND4Bit_1/AND2IN_0/NOT_0/w_n7_n3# 0.03fF
C673 OR3IN_1/vin3 OR2IN_1/vin2 0.06fF
C674 vinSel0 Decoder_0/AND4Bit_0/AND2IN_1/NAND2IN_0/w_n16_n4# 0.10fF
C675 OR2IN_0/vin2 AdderSubtractor_0/fullAdder_0/XOR2IN_1/vin1 0.26fF
C676 OR3IN_2/NOT_0/in OR3IN_2/NOT_0/w_n7_n3# 0.07fF
C677 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_1/w_n16_n4# AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_3/vin1 0.08fF
C678 vdd OR3IN_1/vin1 0.15fF
C679 Comparator_0/NOT_5/out Comparator_0/AND5IN_0/NOT_0/in 0.06fF
C680 AdderSubtractor_0/fullAdder_1/OR2IN_0/vin2 AdderSubtractor_0/fullAdder_1/OR2IN_0/NOT_0/in 0.08fF
C681 OR3IN_2/vin1 vdd 0.15fF
C682 Enable_1/vouta0 Comparator_0/NOT_4/out 0.13fF
C683 AdderSubtractor_0/fullAdder_3/AND2IN_1/NOT_0/w_n7_n3# AdderSubtractor_0/fullAdder_3/AND2IN_1/NOT_0/in 0.07fF
C684 vdd Decoder_0/NOT_1/out 0.06fF
C685 OR2IN_0/NOT_0/w_n7_n3# OR2IN_0/vout 0.03fF
C686 Enable_0/voutb1 Enable_0/vouta2 0.06fF
C687 Enable_0/AND4Bit_1/AND2IN_1/NAND2IN_0/w_n16_n4# vdd 0.11fF
C688 Decoder_0/AND4Bit_0/AND2IN_3/NOT_0/in Decoder_0/AND4Bit_0/AND2IN_3/NOT_0/w_n7_n3# 0.07fF
C689 Enable_2/AND4Bit_0/AND2IN_0/NOT_0/w_n7_n3# vdd 0.06fF
C690 Enable_1/vouta0 Enable_1/vouta3 0.06fF
C691 AND4Bit_0/AND2IN_2/NOT_0/in vdd 0.08fF
C692 Enable_1/AND4Bit_0/AND2IN_0/NAND2IN_0/w_n16_n4# vdd 0.11fF
C693 vdd Decoder_0/AND4Bit_0/AND2IN_0/NOT_0/w_n7_n3# 0.06fF
C694 AdderSubtractor_0/XOR2IN_2/NAND2IN_2/w_n16_n4# AdderSubtractor_0/XOR2IN_2/NAND2IN_2/vin2 0.10fF
C695 Comparator_0/AND2IN_3/NOT_0/w_n7_n3# OR3IN_1/vin2 0.03fF
C696 Comparator_0/AND2IN_1/NOT_0/w_n7_n3# vdd 0.06fF
C697 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_3/w_n16_n4# OR2IN_1/vin1 0.08fF
C698 AND4Bit_0/AND2IN_1/NOT_0/w_n7_n3# vdd 0.06fF
C699 AdderSubtractor_0/XOR2IN_0/NAND2IN_3/w_n16_n4# vdd 0.11fF
C700 OR3IN_1/vin2 OR2IN_1/vin1 0.07fF
C701 Enable_1/vouta3 Comparator_0/XOR2IN_3/NAND2IN_1/w_n16_n4# 0.10fF
C702 vout2 gnd 0.07fF
C703 AdderSubtractor_0/fullAdder_3/AND2IN_0/NOT_0/in AdderSubtractor_0/fullAdder_3/AND2IN_0/NAND2IN_0/w_n16_n4# 0.08fF
C704 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_3/vin2 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_3/w_n16_n4# 0.10fF
C705 Decoder_0/AND4Bit_0/AND2IN_2/NOT_0/in vinSel1 0.06fF
C706 AdderSubtractor_0/XOR2IN_2/NAND2IN_2/w_n16_n4# vdd 0.11fF
C707 Enable_0/AND4Bit_0/AND2IN_0/NAND2IN_0/w_n16_n4# Enable_0/AND4Bit_0/AND2IN_0/NOT_0/in 0.08fF
C708 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_0/w_n16_n4# AdderSubtractor_0/XOR2IN_3/vout 0.10fF
C709 Comparator_0/AND4IN_0/NOT_0/w_n7_n3# Comparator_0/AND4IN_0/vout 0.03fF
C710 gnd AdderSubtractor_0/fullAdder_0/XOR2IN_1/vin1 0.52fF
C711 Enable_2/AND4Bit_1/AND2IN_3/NOT_0/w_n7_n3# Enable_2/AND4Bit_1/AND2IN_3/NOT_0/in 0.07fF
C712 Enable_1/AND4Bit_1/AND2IN_3/NAND2IN_0/w_n16_n4# vdd 0.11fF
C713 Enable_0/voutb2 AdderSubtractor_0/XOR2IN_2/NAND2IN_0/w_n16_n4# 0.10fF
C714 Enable_1/AND4Bit_1/AND2IN_0/NOT_0/w_n7_n3# Enable_1/AND4Bit_1/AND2IN_0/NOT_0/in 0.07fF
C715 Enable_1/voutb2 Comparator_0/NOT_3/out 0.06fF
C716 OR3IN_2/vin2 OR2IN_1/vin1 0.07fF
C717 Comparator_0/AND2IN_3/NAND2IN_0/w_n16_n4# Comparator_0/AND2IN_3/NOT_0/in 0.08fF
C718 AND4Bit_0/AND2IN_1/NAND2IN_0/w_n16_n4# Enable_2/voutb1 0.10fF
C719 Comparator_0/AND4IN_1/w_n14_n10# Comparator_0/NOT_4/out 0.15fF
C720 AdderSubtractor_0/fullAdder_1/vcin vdd 0.12fF
C721 Enable_1/vinEn Enable_1/AND4Bit_0/AND2IN_2/NOT_0/in 0.06fF
C722 vina1 Enable_1/AND4Bit_0/AND2IN_1/NAND2IN_0/w_n16_n4# 0.10fF
C723 Comparator_0/XOR2IN_3/NAND2IN_2/vin2 gnd 0.19fF
C724 Comparator_0/AND2IN_2/NOT_0/w_n7_n3# OR3IN_2/vin2 0.03fF
C725 OR3IN_1/NOT_0/in OR3IN_1/vin3 0.09fF
C726 Comparator_0/AND2IN_3/NOT_0/in gnd 0.05fF
C727 AdderSubtractor_0/XOR2IN_0/NAND2IN_3/w_n16_n4# AdderSubtractor_0/XOR2IN_0/vout 0.08fF
C728 AdderSubtractor_0/fullAdder_1/vcin AdderSubtractor_0/fullAdder_1/OR2IN_0/vin2 0.06fF
C729 vdd Enable_0/vouta1 0.32fF
C730 Comparator_0/XOR2IN_0/NAND2IN_1/w_n16_n4# Comparator_0/XOR2IN_0/NAND2IN_2/vin2 0.10fF
C731 vdd AdderSubtractor_0/fullAdder_0/AND2IN_1/NOT_0/in 0.08fF
C732 AND4Bit_0/AND2IN_0/NOT_0/in Enable_2/voutb0 0.06fF
C733 AdderSubtractor_0/fullAdder_1/XOR2IN_1/vin1 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_3/w_n16_n4# 0.08fF
C734 Comparator_0/NOT_3/out Comparator_0/NOT_4/out 0.13fF
C735 gnd Comparator_0/OR4IN_0/vin3 0.19fF
C736 Comparator_0/AND4IN_0/NOT_0/in gnd 0.03fF
C737 AdderSubtractor_0/XOR2IN_0/NAND2IN_0/w_n16_n4# vdd 0.11fF
C738 Comparator_0/AND5IN_0/w_n26_1# Comparator_0/NOT_4/out 0.12fF
C739 OR3IN_0/vin3 OR3IN_0/NOT_0/in 0.09fF
C740 Enable_1/vinEn Enable_1/AND4Bit_1/AND2IN_1/NOT_0/in 0.06fF
C741 Comparator_0/NOT_6/out gnd 0.39fF
C742 vina0 vina3 0.19fF
C743 Comparator_0/AND2IN_2/NOT_0/in gnd 0.05fF
C744 AdderSubtractor_0/XOR2IN_1/NAND2IN_2/vin2 vdd 0.08fF
C745 gnd vina3 0.19fF
C746 Comparator_0/XOR2IN_3/NAND2IN_3/w_n16_n4# vdd 0.11fF
C747 AdderSubtractor_0/XOR2IN_1/NAND2IN_1/w_n16_n4# AdderSubtractor_0/XOR2IN_1/NAND2IN_2/vin2 0.10fF
C748 Enable_1/vouta3 Comparator_0/NOT_3/out 0.06fF
C749 AND4Bit_0/AND2IN_2/NAND2IN_0/w_n16_n4# Enable_2/voutb2 0.10fF
C750 Enable_1/voutb0 Enable_1/vouta1 0.06fF
C751 Comparator_0/XOR2IN_2/NAND2IN_2/w_n16_n4# Comparator_0/XOR2IN_2/NAND2IN_2/vin2 0.10fF
C752 Comparator_0/NOT_7/in gnd 0.01fF
C753 vina3 Enable_2/AND4Bit_0/AND2IN_3/NAND2IN_0/w_n16_n4# 0.10fF
C754 Enable_2/AND4Bit_0/AND2IN_1/NOT_0/w_n7_n3# Enable_2/vouta1 0.03fF
C755 gnd Enable_2/AND4Bit_0/AND2IN_1/NOT_0/in 0.05fF
C756 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_1/vcin 0.39fF
C757 gnd Enable_1/AND4Bit_0/AND2IN_0/NOT_0/in 0.05fF
C758 OR2IN_0/vout vdd 0.12fF
C759 vina0 vinb2 0.19fF
C760 Comparator_0/XOR2IN_2/NAND2IN_3/vin2 gnd 0.06fF
C761 gnd vinb2 0.19fF
C762 Enable_2/AND4Bit_0/AND2IN_2/NOT_0/in vdd 0.08fF
C763 AdderSubtractor_0/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/XOR2IN_1/NAND2IN_3/vin2 0.06fF
C764 AdderSubtractor_0/fullAdder_2/vcin vdd 0.12fF
C765 Comparator_0/AND3IN_0/NOT_0/w_n7_n3# vdd 0.06fF
C766 OR2IN_1/w_n19_n9# vdd 0.09fF
C767 AdderSubtractor_0/XOR2IN_0/NAND2IN_3/vin2 AdderSubtractor_0/XOR2IN_0/NAND2IN_2/w_n16_n4# 0.08fF
C768 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_0/w_n16_n4# 0.08fF
C769 gnd AdderSubtractor_0/fullAdder_2/XOR2IN_1/vin1 0.52fF
C770 OR3IN_0/vin3 vdd 0.19fF
C771 AdderSubtractor_0/fullAdder_0/AND2IN_0/NOT_0/in vdd 0.08fF
C772 OR2IN_0/vout Enable_0/AND4Bit_0/AND2IN_3/NOT_0/in 0.06fF
C773 Enable_0/voutb0 AdderSubtractor_0/XOR2IN_0/NAND2IN_1/w_n16_n4# 0.10fF
C774 Comparator_0/NOT_5/w_n7_n3# vdd 0.06fF
C775 Decoder_0/AND4Bit_0/AND2IN_2/NAND2IN_0/w_n16_n4# Decoder_0/AND4Bit_0/AND2IN_2/NOT_0/in 0.08fF
C776 Enable_2/AND4Bit_1/AND2IN_1/NOT_0/in vdd 0.08fF
C777 OR2IN_0/vin2 OR2IN_0/vin1 0.11fF
C778 Enable_1/AND4Bit_1/AND2IN_3/NOT_0/w_n7_n3# Enable_1/AND4Bit_1/AND2IN_3/NOT_0/in 0.07fF
C779 Enable_0/AND4Bit_1/AND2IN_0/NOT_0/w_n7_n3# Enable_0/AND4Bit_1/AND2IN_0/NOT_0/in 0.07fF
C780 AND4Bit_0/AND2IN_2/NOT_0/w_n7_n3# vdd 0.06fF
C781 Enable_1/vouta0 vdd 0.32fF
C782 OR2IN_0/vin2 AdderSubtractor_0/XOR2IN_1/NAND2IN_0/w_n16_n4# 0.10fF
C783 vinb2 Enable_2/AND4Bit_1/AND2IN_2/NAND2IN_0/w_n16_n4# 0.10fF
C784 Decoder_0/AND4Bit_0/AND2IN_3/NAND2IN_0/w_n16_n4# vdd 0.11fF
C785 vina2 vinb1 0.19fF
C786 vina1 vinb0 0.19fF
C787 Enable_1/voutb1 Enable_1/vouta2 0.06fF
C788 Enable_1/vouta1 Enable_1/voutb2 0.06fF
C789 OR3IN_0/vin3 AND4Bit_0/AND2IN_0/NOT_0/w_n7_n3# 0.03fF
C790 OR2IN_0/vout Enable_0/AND4Bit_1/AND2IN_2/NOT_0/in 0.06fF
C791 Comparator_0/NOT_7/out Comparator_0/NOT_6/in 0.06fF
C792 Comparator_0/AND2IN_2/NAND2IN_0/w_n16_n4# vdd 0.11fF
C793 gnd AdderSubtractor_0/XOR2IN_1/NAND2IN_3/vin1 0.13fF
C794 Enable_0/AND4Bit_0/AND2IN_2/NAND2IN_0/w_n16_n4# OR2IN_0/vout 0.10fF
C795 Comparator_0/XOR2IN_3/NAND2IN_1/w_n16_n4# vdd 0.11fF
C796 Comparator_0/XOR2IN_1/NAND2IN_1/w_n16_n4# Comparator_0/XOR2IN_1/NAND2IN_2/vin2 0.10fF
C797 Comparator_0/NOT_2/w_n7_n3# Comparator_0/NOT_2/out 0.03fF
C798 AdderSubtractor_0/XOR2IN_0/vout AdderSubtractor_0/fullAdder_0/AND2IN_0/NOT_0/in 0.06fF
C799 Enable_1/vouta1 Comparator_0/NOT_4/out 0.06fF
C800 AdderSubtractor_0/fullAdder_1/XOR2IN_1/vin1 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_3/vin2 0.06fF
C801 Enable_0/vouta0 vdd 0.32fF
C802 Decoder_0/AND4Bit_0/AND2IN_3/NOT_0/w_n7_n3# Enable_2/vinEn 0.03fF
C803 Comparator_0/NOT_6/in vdd 0.19fF
C804 OR3IN_2/w_n19_n9# OR3IN_2/vin1 0.16fF
C805 Enable_1/vouta1 Comparator_0/XOR2IN_1/NAND2IN_0/w_n16_n4# 0.10fF
C806 gnd Enable_2/AND4Bit_1/AND2IN_0/NOT_0/in 0.05fF
C807 Comparator_0/OR4IN_0/NOT_0/w_n7_n3# vdd 0.06fF
C808 Decoder_0/AND4Bit_0/AND2IN_2/NOT_0/w_n7_n3# Enable_1/vinEn 0.03fF
C809 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_3/w_n16_n4# vdd 0.11fF
C810 Enable_1/vouta1 Enable_1/vouta3 0.06fF
C811 Comparator_0/XOR2IN_3/NAND2IN_3/vin2 vdd 0.08fF
C812 Comparator_0/XOR2IN_1/NAND2IN_2/vin2 Comparator_0/XOR2IN_1/NAND2IN_3/vin2 0.06fF
C813 Comparator_0/AND3IN_0/NOT_0/in Comparator_0/NOT_5/out 0.06fF
C814 AdderSubtractor_0/fullAdder_2/vcin Enable_0/vouta2 0.06fF
C815 OR3IN_1/vin2 vdd 0.06fF
C816 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_1/w_n16_n4# AdderSubtractor_0/fullAdder_1/XOR2IN_1/vin1 0.10fF
C817 gnd OR2IN_0/vin1 0.19fF
C818 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_3/vin2 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_3/w_n16_n4# 0.10fF
C819 OR3IN_0/vin2 gnd 0.46fF
C820 Enable_1/AND4Bit_1/AND2IN_0/NOT_0/w_n7_n3# vdd 0.06fF
C821 Enable_0/AND4Bit_0/AND2IN_2/NOT_0/in vdd 0.08fF
C822 Comparator_0/AND4IN_1/w_n14_n10# vdd 0.25fF
C823 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_3/w_n16_n4# AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_3/vin1 0.10fF
C824 gnd Enable_2/vouta0 0.14fF
C825 Comparator_0/AND4IN_0/vout vdd 0.12fF
C826 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_2/w_n16_n4# AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_3/vin2 0.08fF
C827 Comparator_0/NOT_0/w_n7_n3# vdd 0.06fF
C828 gnd AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_2/vin2 0.19fF
C829 OR3IN_2/NOT_0/in OR3IN_2/vin3 0.09fF
C830 Enable_0/vouta0 AdderSubtractor_0/XOR2IN_0/vout 0.27fF
C831 OR3IN_2/vin2 vdd 0.10fF
C832 gnd AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_2/vin2 0.19fF
C833 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_3/w_n16_n4# AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_3/vin1 0.10fF
C834 AND4Bit_0/AND2IN_3/NOT_0/in vdd 0.08fF
C835 Decoder_0/NOT_0/w_n7_n3# vdd 0.06fF
C836 Comparator_0/NOT_3/out vdd 0.06fF
C837 OR3IN_2/vin1 OR3IN_1/vin1 1.64fF
C838 Enable_2/voutb0 vdd 0.19fF
C839 Comparator_0/AND5IN_0/w_n26_1# vdd 0.34fF
C840 AdderSubtractor_0/XOR2IN_2/NAND2IN_2/vin2 AdderSubtractor_0/XOR2IN_2/NAND2IN_3/vin1 0.06fF
C841 Enable_0/AND4Bit_1/AND2IN_1/NOT_0/in vdd 0.08fF
C842 Enable_0/AND4Bit_1/AND2IN_3/NOT_0/w_n7_n3# Enable_0/AND4Bit_1/AND2IN_3/NOT_0/in 0.07fF
C843 Enable_2/vouta1 vdd 0.19fF
C844 Enable_0/voutb0 Enable_0/vouta3 0.46fF
C845 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_2/w_n16_n4# 0.10fF
C846 Enable_0/AND4Bit_1/AND2IN_2/NAND2IN_0/w_n16_n4# vinb2 0.10fF
C847 vdd AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_3/w_n16_n4# 0.11fF
C848 Comparator_0/NOT_5/in Comparator_0/NOT_6/out 0.06fF
C849 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_3/w_n16_n4# vdd 0.11fF
C850 Enable_0/AND4Bit_0/AND2IN_0/NAND2IN_0/w_n16_n4# vdd 0.11fF
C851 AdderSubtractor_0/XOR2IN_2/NAND2IN_3/vin1 vdd 0.43fF
C852 Decoder_0/AND4Bit_0/AND2IN_0/NAND2IN_0/w_n16_n4# Decoder_0/NOT_0/out 0.10fF
C853 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_2/vin2 vdd 0.15fF
C854 AdderSubtractor_0/fullAdder_1/vcin AdderSubtractor_0/fullAdder_1/AND2IN_1/NAND2IN_0/w_n16_n4# 0.10fF
C855 Comparator_0/NOT_2/out Comparator_0/AND4IN_1/NOT_0/in 0.06fF
C856 Decoder_0/AND4Bit_0/AND2IN_1/NAND2IN_0/w_n16_n4# Decoder_0/AND4Bit_0/AND2IN_1/NOT_0/in 0.08fF
C857 Enable_0/AND4Bit_0/AND2IN_2/NAND2IN_0/w_n16_n4# Enable_0/AND4Bit_0/AND2IN_2/NOT_0/in 0.08fF
C858 Decoder_0/AND4Bit_0/AND2IN_0/NOT_0/in Decoder_0/AND4Bit_0/AND2IN_0/NAND2IN_0/w_n16_n4# 0.08fF
C859 vina2 vina3 1.52fF
C860 Enable_1/vinEn Comparator_0/AND2IN_3/NAND2IN_0/w_n16_n4# 0.10fF
C861 Enable_1/voutb3 Comparator_0/XOR2IN_3/NAND2IN_2/w_n16_n4# 0.10fF
C862 vina0 Enable_1/vinEn 0.13fF
C863 Comparator_0/NOT_6/w_n7_n3# Comparator_0/NOT_6/out 0.03fF
C864 AdderSubtractor_0/XOR2IN_1/vout AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_2/vin2 0.39fF
C865 gnd Enable_0/AND4Bit_1/AND2IN_0/NOT_0/in 0.05fF
C866 AdderSubtractor_0/XOR2IN_2/NAND2IN_0/w_n16_n4# AdderSubtractor_0/XOR2IN_2/NAND2IN_2/vin2 0.08fF
C867 vinb0 Enable_2/vinEn 0.19fF
C868 vinSel0 Decoder_0/NOT_0/out 0.06fF
C869 Enable_1/vinEn gnd 1.04fF
C870 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_1/w_n16_n4# 0.10fF
C871 Enable_1/vouta0 Comparator_0/NOT_1/out 0.06fF
C872 Enable_2/vouta2 Enable_2/voutb0 0.06fF
C873 Enable_2/vinEn Enable_2/AND4Bit_0/AND2IN_2/NAND2IN_0/w_n16_n4# 0.10fF
C874 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_3/vin2 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_3/w_n16_n4# 0.10fF
C875 AdderSubtractor_0/XOR2IN_2/vout AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_2/vin2 0.39fF
C876 OR3IN_1/vin3 vdd 0.26fF
C877 AdderSubtractor_0/fullAdder_2/vcin AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_0/w_n16_n4# 0.10fF
C878 vina2 vinb2 0.19fF
C879 AdderSubtractor_0/XOR2IN_2/NAND2IN_0/w_n16_n4# vdd 0.11fF
C880 Enable_2/AND4Bit_1/AND2IN_1/NAND2IN_0/w_n16_n4# Enable_2/AND4Bit_1/AND2IN_1/NOT_0/in 0.08fF
C881 Comparator_0/OR4IN_0/vin2 gnd 0.19fF
C882 Comparator_0/XOR2IN_2/NAND2IN_2/vin2 Comparator_0/XOR2IN_2/NAND2IN_3/vin1 0.06fF
C883 vout1 gnd 0.07fF
C884 Enable_1/AND4Bit_0/AND2IN_2/NOT_0/w_n7_n3# vdd 0.06fF
C885 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_3/w_n16_n4# AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_3/vin1 0.10fF
C886 vdd AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_1/w_n16_n4# 0.11fF
C887 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_1/w_n16_n4# vdd 0.11fF
C888 Enable_0/voutb0 vdd 0.32fF
C889 Enable_1/vouta0 Enable_1/voutb1 0.06fF
C890 Comparator_0/AND2IN_3/NOT_0/w_n7_n3# Comparator_0/AND2IN_3/NOT_0/in 0.07fF
C891 Enable_1/vouta1 vdd 0.32fF
C892 gnd AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_3/vin1 0.06fF
C893 AdderSubtractor_0/fullAdder_2/vcin AdderSubtractor_0/fullAdder_2/AND2IN_1/NAND2IN_0/w_n16_n4# 0.10fF
C894 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_0/w_n16_n4# AdderSubtractor_0/fullAdder_0/XOR2IN_1/vin1 0.10fF
C895 AdderSubtractor_0/fullAdder_3/OR2IN_0/vin1 AdderSubtractor_0/fullAdder_3/OR2IN_0/w_n19_n9# 0.16fF
C896 gnd AND4Bit_0/AND2IN_1/NOT_0/in 0.05fF
C897 Enable_1/AND4Bit_1/AND2IN_1/NOT_0/w_n7_n3# vdd 0.06fF
C898 OR2IN_1/NOT_0/in OR2IN_1/NOT_0/w_n7_n3# 0.07fF
C899 vdd AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_3/vin2 0.08fF
C900 Comparator_0/AND4IN_0/NOT_0/w_n7_n3# Comparator_0/AND4IN_0/NOT_0/in 0.07fF
C901 AdderSubtractor_0/XOR2IN_3/vout AdderSubtractor_0/XOR2IN_3/NAND2IN_3/w_n16_n4# 0.08fF
C902 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_3/vin2 vdd 0.08fF
C903 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_1/w_n16_n4# AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_2/vin2 0.10fF
C904 Comparator_0/XOR2IN_2/NAND2IN_0/w_n16_n4# Comparator_0/XOR2IN_2/NAND2IN_2/vin2 0.08fF
C905 AdderSubtractor_0/fullAdder_0/AND2IN_1/NAND2IN_0/w_n16_n4# vdd 0.14fF
C906 OR2IN_0/vout Enable_0/AND4Bit_1/AND2IN_1/NAND2IN_0/w_n16_n4# 0.10fF
C907 Comparator_0/AND4IN_0/NOT_0/in Comparator_0/NOT_4/out 0.06fF
C908 Comparator_0/AND2IN_2/NOT_0/w_n7_n3# Comparator_0/AND2IN_2/NOT_0/in 0.07fF
C909 OR3IN_0/vin3 OR3IN_1/vin1 0.07fF
C910 Enable_1/vouta0 Enable_1/vouta2 0.06fF
C911 gnd vcout 0.07fF
C912 AdderSubtractor_0/fullAdder_1/vcin Enable_0/vouta1 0.06fF
C913 vdd AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_1/w_n16_n4# 0.11fF
C914 gnd Enable_1/AND4Bit_0/AND2IN_3/NOT_0/in 0.05fF
C915 gnd Comparator_0/OR4IN_0/vout 0.14fF
C916 OR3IN_0/vin3 OR3IN_2/vin1 0.07fF
C917 vdd AdderSubtractor_0/fullAdder_0/AND2IN_0/NOT_0/w_n7_n3# 0.09fF
C918 gnd Comparator_0/AND4IN_1/NOT_0/in 0.03fF
C919 Enable_0/vouta3 AdderSubtractor_0/fullAdder_3/AND2IN_0/NAND2IN_0/w_n16_n4# 0.10fF
C920 AND4Bit_0/AND2IN_3/NOT_0/in AND4Bit_0/AND2IN_3/NAND2IN_0/w_n16_n4# 0.08fF
C921 AdderSubtractor_0/fullAdder_3/vcin AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_0/w_n16_n4# 0.10fF
C922 Enable_2/vinEn Enable_2/AND4Bit_0/AND2IN_0/NAND2IN_0/w_n16_n4# 0.10fF
C923 Enable_1/vouta3 Comparator_0/NOT_6/out 0.06fF
C924 AdderSubtractor_0/XOR2IN_1/NAND2IN_2/w_n16_n4# vdd 0.11fF
C925 Enable_1/AND4Bit_1/AND2IN_1/NAND2IN_0/w_n16_n4# Enable_1/AND4Bit_1/AND2IN_1/NOT_0/in 0.08fF
C926 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_1/w_n16_n4# AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_3/vin1 0.08fF
C927 OR3IN_0/vin1 vdd 0.24fF
C928 gnd Enable_1/AND4Bit_1/AND2IN_2/NOT_0/in 0.05fF
C929 Comparator_0/AND5IN_0/NOT_0/in gnd 0.03fF
C930 Enable_0/voutb0 Enable_0/vouta2 0.06fF
C931 Enable_0/vouta2 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_1/w_n16_n4# 0.10fF
C932 Enable_1/voutb1 Comparator_0/NOT_3/out 0.06fF
C933 Comparator_0/XOR2IN_0/NAND2IN_0/w_n16_n4# Comparator_0/XOR2IN_0/NAND2IN_2/vin2 0.08fF
C934 Enable_2/AND4Bit_0/AND2IN_1/NOT_0/w_n7_n3# Enable_2/AND4Bit_0/AND2IN_1/NOT_0/in 0.07fF
C935 Comparator_0/AND2IN_1/NAND2IN_0/w_n16_n4# vdd 0.11fF
C936 OR3IN_2/w_n19_n9# OR3IN_2/vin2 0.12fF
C937 Enable_1/AND4Bit_1/AND2IN_3/NOT_0/in vdd 0.08fF
C938 AND4Bit_0/AND2IN_2/NOT_0/w_n7_n3# AND4Bit_0/AND2IN_2/NOT_0/in 0.07fF
C939 Comparator_0/XOR2IN_2/NAND2IN_2/vin2 gnd 0.19fF
C940 vout1 OR3IN_1/NOT_0/w_n7_n3# 0.03fF
C941 AdderSubtractor_0/fullAdder_0/OR2IN_0/NOT_0/in AdderSubtractor_0/fullAdder_0/OR2IN_0/w_n19_n9# 0.05fF
C942 Enable_2/vinEn Enable_2/AND4Bit_1/AND2IN_3/NAND2IN_0/w_n16_n4# 0.10fF
C943 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_1/w_n16_n4# AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_2/vin2 0.10fF
C944 Comparator_0/XOR2IN_0/NAND2IN_1/w_n16_n4# vdd 0.11fF
C945 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_1/w_n16_n4# 0.10fF
C946 vinb3 Enable_1/AND4Bit_1/AND2IN_3/NAND2IN_0/w_n16_n4# 0.10fF
C947 AdderSubtractor_0/XOR2IN_1/NAND2IN_2/w_n16_n4# AdderSubtractor_0/XOR2IN_1/NAND2IN_3/vin2 0.08fF
C948 OR2IN_0/vin2 AdderSubtractor_0/XOR2IN_0/NAND2IN_2/w_n16_n4# 0.10fF
C949 Enable_0/AND4Bit_0/AND2IN_1/NOT_0/in Enable_0/AND4Bit_0/AND2IN_1/NOT_0/w_n7_n3# 0.07fF
C950 OR3IN_1/vin2 OR3IN_1/vin1 0.14fF
C951 AdderSubtractor_0/XOR2IN_0/NAND2IN_2/vin2 AdderSubtractor_0/XOR2IN_0/NAND2IN_2/w_n16_n4# 0.10fF
C952 Comparator_0/AND3IN_0/w_n14_n10# vdd 0.19fF
C953 Decoder_0/AND4Bit_0/AND2IN_2/NAND2IN_0/w_n16_n4# vdd 0.11fF
C954 OR3IN_1/vin2 OR3IN_2/vin1 0.07fF
C955 AND4Bit_0/AND2IN_2/NAND2IN_0/w_n16_n4# vdd 0.11fF
C956 Comparator_0/XOR2IN_2/NAND2IN_3/w_n16_n4# vdd 0.11fF
C957 Enable_1/vouta2 Comparator_0/NOT_3/out 0.06fF
C958 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_3/vin2 0.06fF
C959 vina1 Enable_2/vinEn 0.19fF
C960 Enable_1/AND4Bit_0/AND2IN_3/NAND2IN_0/w_n16_n4# vdd 0.11fF
C961 Comparator_0/AND2IN_0/NOT_0/w_n7_n3# vdd 0.06fF
C962 AdderSubtractor_0/XOR2IN_3/NAND2IN_3/vin2 AdderSubtractor_0/XOR2IN_3/NAND2IN_3/w_n16_n4# 0.10fF
C963 OR2IN_0/w_n19_n9# OR2IN_0/vin2 0.12fF
C964 AdderSubtractor_0/fullAdder_3/OR2IN_0/NOT_0/w_n7_n3# AdderSubtractor_0/fullAdder_3/OR2IN_0/NOT_0/in 0.07fF
C965 AND4Bit_0/AND2IN_1/NAND2IN_0/w_n16_n4# Enable_2/vouta1 0.10fF
C966 OR2IN_0/vin2 Decoder_0/AND4Bit_0/AND2IN_1/NOT_0/w_n7_n3# 0.03fF
C967 OR3IN_2/vin2 OR3IN_2/vin1 0.14fF
C968 AdderSubtractor_0/XOR2IN_3/vout AdderSubtractor_0/XOR2IN_3/NAND2IN_3/vin2 0.06fF
C969 Comparator_0/XOR2IN_1/NAND2IN_3/vin2 gnd 0.06fF
C970 AdderSubtractor_0/XOR2IN_0/NAND2IN_2/vin2 AdderSubtractor_0/XOR2IN_0/NAND2IN_3/vin1 0.06fF
C971 AdderSubtractor_0/fullAdder_3/AND2IN_0/NAND2IN_0/w_n16_n4# vdd 0.11fF
C972 Enable_1/vouta1 Comparator_0/NOT_1/out 0.06fF
C973 Enable_1/vinEn vina2 0.13fF
C974 Enable_1/AND4Bit_1/AND2IN_2/NAND2IN_0/w_n16_n4# vdd 0.11fF
C975 Enable_1/vinEn Enable_1/AND4Bit_1/AND2IN_0/NAND2IN_0/w_n16_n4# 0.10fF
C976 OR2IN_0/vout vinb3 0.06fF
C977 vout2 vdd 0.24fF
C978 OR3IN_0/vin2 OR2IN_1/vin1 0.07fF
C979 Enable_1/vinEn Enable_1/AND4Bit_0/AND2IN_1/NOT_0/in 0.06fF
C980 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_0/w_n16_n4# vdd 0.11fF
C981 AdderSubtractor_0/fullAdder_0/XOR2IN_1/vin1 vdd 0.21fF
C982 AdderSubtractor_0/fullAdder_2/XOR2IN_1/vin1 AdderSubtractor_0/fullAdder_2/AND2IN_1/NOT_0/in 0.06fF
C983 Enable_0/AND4Bit_1/AND2IN_1/NAND2IN_0/w_n16_n4# Enable_0/AND4Bit_1/AND2IN_1/NOT_0/in 0.08fF
C984 gnd Decoder_0/NOT_0/out 0.26fF
C985 Comparator_0/NOT_7/out Comparator_0/NOT_6/out 0.06fF
C986 Comparator_0/XOR2IN_0/NAND2IN_3/vin2 Comparator_0/XOR2IN_0/NAND2IN_3/w_n16_n4# 0.10fF
C987 AdderSubtractor_0/XOR2IN_1/vout AdderSubtractor_0/fullAdder_1/AND2IN_0/NAND2IN_0/w_n16_n4# 0.10fF
C988 AdderSubtractor_0/fullAdder_3/AND2IN_1/NOT_0/w_n7_n3# vdd 0.06fF
C989 AdderSubtractor_0/fullAdder_3/vcin AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_2/w_n16_n4# 0.10fF
C990 Comparator_0/NOT_5/out Comparator_0/NOT_0/out 0.06fF
C991 OR2IN_1/vin2 vcout 0.06fF
C992 AdderSubtractor_0/fullAdder_1/AND2IN_1/NOT_0/w_n7_n3# AdderSubtractor_0/fullAdder_1/OR2IN_0/vin1 0.03fF
C993 Enable_1/AND4Bit_0/AND2IN_1/NOT_0/w_n7_n3# Enable_1/AND4Bit_0/AND2IN_1/NOT_0/in 0.07fF
C994 AND4Bit_0/AND2IN_2/NAND2IN_0/w_n16_n4# Enable_2/vouta2 0.10fF
C995 Comparator_0/XOR2IN_3/NAND2IN_2/vin2 vdd 0.08fF
C996 Comparator_0/XOR2IN_1/NAND2IN_2/w_n16_n4# Comparator_0/XOR2IN_1/NAND2IN_3/vin2 0.08fF
C997 Comparator_0/NOT_5/out Comparator_0/NOT_2/out 0.13fF
C998 Enable_0/voutb0 Enable_0/voutb1 1.49fF
C999 vina0 vinb0 0.19fF
C1000 AdderSubtractor_0/fullAdder_0/OR2IN_0/vin2 AdderSubtractor_0/fullAdder_0/AND2IN_0/NOT_0/w_n7_n3# 0.03fF
C1001 Comparator_0/AND2IN_3/NOT_0/in vdd 0.08fF
C1002 AdderSubtractor_0/XOR2IN_2/vout AdderSubtractor_0/fullAdder_2/AND2IN_0/NAND2IN_0/w_n16_n4# 0.10fF
C1003 Enable_1/vouta1 Enable_1/voutb1 0.06fF
C1004 gnd vinb0 0.19fF
C1005 Comparator_0/OR4IN_0/w_n19_n9# vdd 0.11fF
C1006 gnd Decoder_0/AND4Bit_0/AND2IN_0/NOT_0/in 0.05fF
C1007 AdderSubtractor_0/fullAdder_2/AND2IN_1/NOT_0/w_n7_n3# AdderSubtractor_0/fullAdder_2/OR2IN_0/vin1 0.03fF
C1008 Comparator_0/AND2IN_1/NOT_0/in gnd 0.05fF
C1009 Comparator_0/OR4IN_0/vin3 vdd 0.20fF
C1010 Comparator_0/AND4IN_0/NOT_0/in vdd 0.26fF
C1011 AdderSubtractor_0/fullAdder_0/OR2IN_0/vin2 AdderSubtractor_0/fullAdder_0/OR2IN_0/NOT_0/in 0.08fF
C1012 Enable_2/AND4Bit_1/AND2IN_3/NOT_0/w_n7_n3# vdd 0.06fF
C1013 Enable_1/voutb1 Enable_1/AND4Bit_1/AND2IN_1/NOT_0/w_n7_n3# 0.03fF
C1014 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_2/w_n16_n4# AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_2/vin2 0.10fF
C1015 gnd AdderSubtractor_0/XOR2IN_0/NAND2IN_3/vin1 0.13fF
C1016 Comparator_0/XOR2IN_2/NAND2IN_1/w_n16_n4# vdd 0.11fF
C1017 Enable_2/AND4Bit_0/AND2IN_1/NAND2IN_0/w_n16_n4# Enable_2/AND4Bit_0/AND2IN_1/NOT_0/in 0.08fF
C1018 Comparator_0/XOR2IN_2/NAND2IN_3/w_n16_n4# Comparator_0/NOT_4/in 0.08fF
C1019 Comparator_0/NOT_6/out vdd 0.12fF
C1020 Comparator_0/AND2IN_2/NOT_0/in vdd 0.08fF
C1021 Enable_0/voutb3 AdderSubtractor_0/XOR2IN_3/NAND2IN_1/w_n16_n4# 0.10fF
C1022 Comparator_0/XOR2IN_0/NAND2IN_0/w_n16_n4# Enable_1/voutb0 0.10fF
C1023 AdderSubtractor_0/XOR2IN_1/NAND2IN_3/w_n16_n4# AdderSubtractor_0/XOR2IN_1/NAND2IN_3/vin1 0.10fF
C1024 Comparator_0/XOR2IN_3/NAND2IN_3/vin2 Comparator_0/XOR2IN_3/NAND2IN_3/w_n16_n4# 0.10fF
C1025 Comparator_0/XOR2IN_3/NAND2IN_0/w_n16_n4# Enable_1/voutb3 0.10fF
C1026 Enable_2/AND4Bit_1/AND2IN_0/NAND2IN_0/w_n16_n4# vdd 0.11fF
C1027 Enable_1/vouta2 Enable_1/AND4Bit_0/AND2IN_2/NOT_0/w_n7_n3# 0.03fF
C1028 Comparator_0/NOT_7/in vdd 0.19fF
C1029 Enable_2/AND4Bit_0/AND2IN_1/NOT_0/in vdd 0.08fF
C1030 Enable_1/AND4Bit_0/AND2IN_0/NOT_0/in vdd 0.08fF
C1031 Comparator_0/XOR2IN_2/NAND2IN_3/vin2 vdd 0.08fF
C1032 Enable_2/AND4Bit_0/AND2IN_3/NOT_0/w_n7_n3# Enable_2/vouta3 0.03fF
C1033 Enable_1/vouta1 Enable_1/vouta2 27.66fF
C1034 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_2/w_n16_n4# vdd 0.11fF
C1035 OR2IN_0/vout Enable_0/AND4Bit_0/AND2IN_2/NOT_0/in 0.06fF
C1036 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_2/w_n16_n4# AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_3/vin2 0.08fF
C1037 vinb1 Enable_2/AND4Bit_1/AND2IN_1/NAND2IN_0/w_n16_n4# 0.10fF
C1038 Enable_1/vinEn Enable_1/AND4Bit_1/AND2IN_0/NOT_0/in 0.06fF
C1039 AND4Bit_0/AND2IN_1/NOT_0/w_n7_n3# OR3IN_1/vin3 0.03fF
C1040 Decoder_0/NOT_0/out Decoder_0/AND4Bit_0/AND2IN_1/NOT_0/in 0.06fF
C1041 AdderSubtractor_0/fullAdder_2/XOR2IN_1/vin1 vdd 0.21fF
C1042 Comparator_0/XOR2IN_3/NAND2IN_3/vin1 gnd 0.13fF
C1043 OR3IN_0/vin3 OR3IN_1/vin2 0.07fF
C1044 Comparator_0/AND3IN_0/w_n14_n10# Comparator_0/NOT_1/out 0.15fF
C1045 Comparator_0/XOR2IN_0/NAND2IN_1/w_n16_n4# Comparator_0/XOR2IN_0/NAND2IN_3/vin1 0.08fF
C1046 AdderSubtractor_0/XOR2IN_1/vout AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_2/w_n16_n4# 0.10fF
C1047 OR2IN_0/vout Enable_0/AND4Bit_1/AND2IN_1/NOT_0/in 0.06fF
C1048 OR3IN_2/vin3 gnd 0.26fF
C1049 vinSel1 Decoder_0/NOT_1/out 0.09fF
C1050 OR3IN_0/vin2 OR3IN_0/NOT_0/in 0.08fF
C1051 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_2/w_n16_n4# vdd 0.11fF
C1052 Enable_0/AND4Bit_0/AND2IN_1/NOT_0/w_n7_n3# vdd 0.06fF
C1053 vdd AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_3/w_n16_n4# 0.11fF
C1054 OR3IN_0/vin3 OR3IN_2/vin2 7.72fF
C1055 AdderSubtractor_0/XOR2IN_2/vout AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_2/w_n16_n4# 0.10fF
C1056 Enable_2/AND4Bit_1/AND2IN_2/NOT_0/w_n7_n3# Enable_2/voutb2 0.03fF
C1057 Enable_0/AND4Bit_0/AND2IN_0/NAND2IN_0/w_n16_n4# OR2IN_0/vout 0.10fF
C1058 Comparator_0/NOT_4/in Comparator_0/NOT_6/out 0.06fF
C1059 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_3/w_n16_n4# vdd 0.11fF
C1060 Enable_2/vinEn vinSel0 0.03fF
C1061 Decoder_0/AND4Bit_0/AND2IN_1/NOT_0/w_n7_n3# Decoder_0/AND4Bit_0/AND2IN_1/NOT_0/in 0.07fF
C1062 AdderSubtractor_0/XOR2IN_1/NAND2IN_3/vin1 vdd 0.43fF
C1063 Comparator_0/XOR2IN_1/NAND2IN_3/w_n16_n4# Comparator_0/XOR2IN_1/NAND2IN_3/vin1 0.10fF
C1064 Comparator_0/AND3IN_0/NOT_0/in gnd 0.06fF
C1065 AdderSubtractor_0/XOR2IN_1/NAND2IN_1/w_n16_n4# AdderSubtractor_0/XOR2IN_1/NAND2IN_3/vin1 0.08fF
C1066 vina0 Enable_2/AND4Bit_0/AND2IN_0/NAND2IN_0/w_n16_n4# 0.10fF
C1067 Enable_0/AND4Bit_1/AND2IN_3/NOT_0/w_n7_n3# vdd 0.06fF
C1068 Enable_2/AND4Bit_1/AND2IN_3/NAND2IN_0/w_n16_n4# Enable_2/AND4Bit_1/AND2IN_3/NOT_0/in 0.08fF
C1069 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_3/vin2 0.06fF
C1070 Enable_1/AND4Bit_0/AND2IN_1/NAND2IN_0/w_n16_n4# Enable_1/AND4Bit_0/AND2IN_1/NOT_0/in 0.08fF
C1071 AdderSubtractor_0/XOR2IN_0/NAND2IN_2/vin2 AdderSubtractor_0/XOR2IN_0/NAND2IN_3/vin2 0.06fF
C1072 Comparator_0/NOT_5/out gnd 0.45fF
C1073 gnd AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_2/vin2 0.19fF
C1074 vdd Decoder_0/AND4Bit_0/AND2IN_1/NAND2IN_0/w_n16_n4# 0.11fF
C1075 Enable_1/vouta0 Comparator_0/AND5IN_0/w_n26_1# 0.12fF
C1076 Comparator_0/XOR2IN_2/NAND2IN_3/vin2 Comparator_0/NOT_4/in 0.06fF
C1077 AdderSubtractor_0/fullAdder_3/OR2IN_0/NOT_0/w_n7_n3# vdd 0.09fF
C1078 Enable_2/AND4Bit_1/AND2IN_0/NOT_0/in vdd 0.08fF
C1079 Enable_0/AND4Bit_1/AND2IN_0/NAND2IN_0/w_n16_n4# vdd 0.11fF
C1080 AdderSubtractor_0/XOR2IN_3/vout OR2IN_0/vin2 0.06fF
C1081 Comparator_0/OR4IN_0/vin1 gnd 0.19fF
C1082 Enable_0/vouta1 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_1/w_n16_n4# 0.10fF
C1083 Decoder_0/AND4Bit_0/AND2IN_3/NOT_0/in gnd 0.05fF
C1084 Enable_0/voutb0 Enable_0/vouta1 0.06fF
C1085 vdd OR2IN_0/vin1 0.19fF
C1086 OR3IN_0/vin2 vdd 0.16fF
C1087 vout3 OR2IN_1/NOT_0/w_n7_n3# 0.03fF
C1088 Comparator_0/AND4IN_1/NOT_0/w_n7_n3# Comparator_0/OR4IN_0/vin3 0.03fF
C1089 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_3/w_n16_n4# vdd 0.11fF
C1090 Enable_0/voutb0 AdderSubtractor_0/XOR2IN_0/NAND2IN_0/w_n16_n4# 0.10fF
C1091 Enable_2/vouta0 vdd 0.19fF
C1092 AdderSubtractor_0/XOR2IN_1/NAND2IN_0/w_n16_n4# vdd 0.11fF
C1093 vdd AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_2/vin2 0.15fF
C1094 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_2/vin2 vdd 0.15fF
C1095 vinb1 Enable_0/AND4Bit_1/AND2IN_1/NAND2IN_0/w_n16_n4# 0.10fF
C1096 Comparator_0/AND3IN_0/w_n14_n10# Enable_1/vouta2 0.15fF
C1097 OR3IN_2/NOT_0/in gnd 0.26fF
C1098 Comparator_0/NOT_6/out Comparator_0/NOT_1/out 0.06fF
C1099 Comparator_0/AND4IN_1/NOT_0/in Comparator_0/NOT_4/out 0.06fF
C1100 OR3IN_2/vin2 OR3IN_1/vin2 7.21fF
C1101 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_1/w_n16_n4# AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_3/vin1 0.08fF
C1102 vina1 Enable_0/AND4Bit_0/AND2IN_1/NAND2IN_0/w_n16_n4# 0.10fF
C1103 vina0 vina1 3.35fF
C1104 Comparator_0/AND4IN_0/NOT_0/in Comparator_0/AND4IN_0/w_n14_n10# 0.25fF
C1105 Comparator_0/OR4IN_0/vin4 Comparator_0/OR4IN_0/w_n19_n9# 0.12fF
C1106 gnd AdderSubtractor_0/XOR2IN_0/NAND2IN_3/vin2 0.06fF
C1107 vina1 gnd 0.19fF
C1108 Comparator_0/OR4IN_0/vin4 Comparator_0/OR4IN_0/vin3 1.01fF
C1109 gnd AdderSubtractor_0/fullAdder_3/OR2IN_0/vin1 0.26fF
C1110 Comparator_0/NOT_6/out Comparator_0/AND4IN_0/w_n14_n10# 0.15fF
C1111 gnd Comparator_0/OR4IN_0/NOT_0/in 0.36fF
C1112 Enable_1/voutb2 Comparator_0/XOR2IN_2/NAND2IN_2/vin2 0.39fF
C1113 AdderSubtractor_0/fullAdder_0/AND2IN_1/NAND2IN_0/w_n16_n4# AdderSubtractor_0/fullAdder_0/AND2IN_1/NOT_0/in 0.08fF
C1114 gnd AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_3/vin1 0.06fF
C1115 Comparator_0/XOR2IN_1/NAND2IN_1/w_n16_n4# Comparator_0/XOR2IN_1/NAND2IN_3/vin1 0.08fF
C1116 Comparator_0/AND5IN_0/NOT_0/in Comparator_0/NOT_4/out 0.06fF
C1117 Decoder_0/AND4Bit_0/AND2IN_2/NAND2IN_0/w_n16_n4# Decoder_0/NOT_1/out 0.10fF
C1118 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_3/vin2 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_2/w_n16_n4# 0.08fF
C1119 Comparator_0/NOR2IN_0/vout Comparator_0/AND2IN_3/NAND2IN_0/w_n16_n4# 0.10fF
C1120 vina2 vinb0 0.19fF
C1121 gnd AdderSubtractor_0/XOR2IN_3/vout 0.28fF
C1122 gnd Enable_2/voutb3 0.14fF
C1123 vout3 OR3IN_2/vin3 0.06fF
C1124 vina2 Enable_2/AND4Bit_0/AND2IN_2/NAND2IN_0/w_n16_n4# 0.10fF
C1125 vinb0 Enable_1/AND4Bit_1/AND2IN_0/NAND2IN_0/w_n16_n4# 0.10fF
C1126 Comparator_0/NOR2IN_0/vout gnd 0.17fF
C1127 Comparator_0/AND5IN_0/w_n26_1# Comparator_0/NOT_3/out 0.12fF
C1128 Enable_1/AND4Bit_1/AND2IN_3/NAND2IN_0/w_n16_n4# Enable_1/AND4Bit_1/AND2IN_3/NOT_0/in 0.08fF
C1129 AND4Bit_0/AND2IN_2/NAND2IN_0/w_n16_n4# AND4Bit_0/AND2IN_2/NOT_0/in 0.08fF
C1130 AdderSubtractor_0/XOR2IN_3/vout AdderSubtractor_0/fullAdder_3/AND2IN_0/NOT_0/in 0.06fF
C1131 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_3/vin2 vdd 0.08fF
C1132 Comparator_0/NOR2IN_0/w_n19_n9# vdd 0.09fF
C1133 gnd AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_2/vin2 0.19fF
C1134 AdderSubtractor_0/fullAdder_1/XOR2IN_1/vin1 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_0/w_n16_n4# 0.10fF
C1135 Decoder_0/NOT_1/w_n7_n3# vinSel0 0.07fF
C1136 OR3IN_2/vin3 OR2IN_1/vin2 7.61fF
C1137 Enable_2/vouta1 Enable_2/voutb0 0.06fF
C1138 Enable_2/AND4Bit_0/AND2IN_0/NAND2IN_0/w_n16_n4# Enable_2/AND4Bit_0/AND2IN_0/NOT_0/in 0.08fF
C1139 Enable_0/AND4Bit_1/AND2IN_0/NOT_0/in vdd 0.08fF
C1140 Enable_1/vouta0 Enable_1/vouta1 28.47fF
C1141 AdderSubtractor_0/fullAdder_3/OR2IN_0/vin2 AdderSubtractor_0/fullAdder_3/OR2IN_0/vin1 0.11fF
C1142 Enable_1/vinEn vdd 0.52fF
C1143 Enable_0/voutb3 OR2IN_0/vin2 0.06fF
C1144 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_3/vin1 0.06fF
C1145 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_1/w_n16_n4# vdd 0.11fF
C1146 AdderSubtractor_0/XOR2IN_1/NAND2IN_2/w_n16_n4# AdderSubtractor_0/XOR2IN_1/NAND2IN_2/vin2 0.10fF
C1147 Comparator_0/NOT_2/w_n7_n3# vdd 0.06fF
C1148 gnd AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_3/vin1 0.06fF
C1149 Enable_0/vouta3 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_0/w_n16_n4# 0.10fF
C1150 gnd AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_3/vin1 0.06fF
C1151 Decoder_0/AND4Bit_0/AND2IN_3/NAND2IN_0/w_n16_n4# vinSel1 0.10fF
C1152 AdderSubtractor_0/fullAdder_3/OR2IN_0/vin2 AdderSubtractor_0/fullAdder_3/OR2IN_0/w_n19_n9# 0.12fF
C1153 Enable_1/vouta2 Comparator_0/XOR2IN_2/NAND2IN_1/w_n16_n4# 0.10fF
C1154 OR3IN_1/vin2 OR3IN_1/vin3 0.14fF
C1155 Enable_1/AND4Bit_0/AND2IN_1/NOT_0/w_n7_n3# vdd 0.06fF
C1156 Enable_1/vouta2 Comparator_0/NOT_6/out 0.06fF
C1157 Comparator_0/OR4IN_0/vin2 vdd 0.22fF
C1158 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_0/w_n16_n4# AdderSubtractor_0/fullAdder_2/XOR2IN_1/vin1 0.10fF
C1159 vout1 vdd 0.24fF
C1160 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_2/w_n16_n4# AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_3/vin2 0.08fF
C1161 OR2IN_0/vout vinb1 0.06fF
C1162 Comparator_0/XOR2IN_0/NAND2IN_0/w_n16_n4# vdd 0.11fF
C1163 AdderSubtractor_0/fullAdder_0/AND2IN_0/NOT_0/in AdderSubtractor_0/fullAdder_0/AND2IN_0/NOT_0/w_n7_n3# 0.07fF
C1164 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_3/vin2 vdd 0.08fF
C1165 Comparator_0/XOR2IN_1/NAND2IN_2/vin2 gnd 0.19fF
C1166 AdderSubtractor_0/XOR2IN_0/NAND2IN_1/w_n16_n4# AdderSubtractor_0/XOR2IN_0/NAND2IN_3/vin1 0.08fF
C1167 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_3/vin1 vdd 0.43fF
C1168 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_3/vin1 0.06fF
C1169 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_3/vin1 0.06fF
C1170 vinb1 vinb3 0.19fF
C1171 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_0/w_n16_n4# AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_2/vin2 0.08fF
C1172 AND4Bit_0/AND2IN_1/NOT_0/in vdd 0.08fF
C1173 AdderSubtractor_0/fullAdder_2/XOR2IN_1/vin1 AdderSubtractor_0/fullAdder_2/AND2IN_1/NAND2IN_0/w_n16_n4# 0.10fF
C1174 Enable_2/vinEn Enable_2/AND4Bit_1/AND2IN_3/NOT_0/in 0.06fF
C1175 Enable_1/vouta1 Comparator_0/AND4IN_1/w_n14_n10# 0.15fF
C1176 Enable_0/AND4Bit_1/AND2IN_2/NOT_0/w_n7_n3# Enable_0/voutb2 0.03fF
C1177 Comparator_0/NOT_5/out Comparator_0/NOT_5/in 0.06fF
C1178 gnd Enable_0/voutb3 0.34fF
C1179 Comparator_0/XOR2IN_1/NAND2IN_3/w_n16_n4# vdd 0.11fF
C1180 OR3IN_2/NOT_0/w_n7_n3# vdd 0.06fF
C1181 gnd AdderSubtractor_0/XOR2IN_3/NAND2IN_3/vin2 0.06fF
C1182 gnd Enable_1/AND4Bit_0/AND2IN_2/NOT_0/in 0.05fF
C1183 Enable_0/AND4Bit_1/AND2IN_3/NAND2IN_0/w_n16_n4# Enable_0/AND4Bit_1/AND2IN_3/NOT_0/in 0.08fF
C1184 Enable_1/vouta1 Comparator_0/NOT_3/out 0.06fF
C1185 AdderSubtractor_0/fullAdder_1/AND2IN_1/NOT_0/w_n7_n3# AdderSubtractor_0/fullAdder_1/AND2IN_1/NOT_0/in 0.07fF
C1186 vina0 Enable_2/vinEn 0.19fF
C1187 Comparator_0/XOR2IN_3/NAND2IN_2/w_n16_n4# vdd 0.11fF
C1188 AdderSubtractor_0/fullAdder_0/XOR2IN_1/vin1 AdderSubtractor_0/fullAdder_0/AND2IN_1/NOT_0/in 0.06fF
C1189 Comparator_0/XOR2IN_1/NAND2IN_2/w_n16_n4# Comparator_0/XOR2IN_1/NAND2IN_2/vin2 0.10fF
C1190 gnd Enable_2/vinEn 0.65fF
C1191 vcout vdd 0.12fF
C1192 Decoder_0/NOT_0/w_n7_n3# vinSel1 0.07fF
C1193 Enable_1/AND4Bit_0/AND2IN_3/NOT_0/in vdd 0.08fF
C1194 Comparator_0/XOR2IN_0/NAND2IN_3/vin2 gnd 0.06fF
C1195 Comparator_0/OR4IN_0/vout vdd 0.08fF
C1196 Comparator_0/NOT_0/out Comparator_0/AND2IN_0/NOT_0/in 0.06fF
C1197 AdderSubtractor_0/fullAdder_2/AND2IN_1/NOT_0/w_n7_n3# AdderSubtractor_0/fullAdder_2/AND2IN_1/NOT_0/in 0.07fF
C1198 Enable_1/AND4Bit_0/AND2IN_0/NAND2IN_0/w_n16_n4# Enable_1/AND4Bit_0/AND2IN_0/NOT_0/in 0.08fF
C1199 Comparator_0/AND4IN_1/NOT_0/in vdd 0.26fF
C1200 Enable_1/vouta0 Comparator_0/XOR2IN_0/NAND2IN_1/w_n16_n4# 0.10fF
C1201 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_0/w_n16_n4# vdd 0.11fF
C1202 Enable_2/vinEn Enable_2/AND4Bit_0/AND2IN_3/NAND2IN_0/w_n16_n4# 0.10fF
C1203 Comparator_0/AND5IN_0/NOT_0/w_n7_n3# Comparator_0/AND5IN_0/NOT_0/in 0.07fF
C1204 Enable_1/voutb3 Comparator_0/NOT_2/out 0.06fF
C1205 gnd Enable_1/AND4Bit_1/AND2IN_1/NOT_0/in 0.05fF
C1206 gnd vinSel0 0.20fF
C1207 Enable_0/voutb1 AdderSubtractor_0/XOR2IN_1/NAND2IN_0/w_n16_n4# 0.10fF
C1208 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_3/w_n16_n4# OR3IN_1/vin1 0.08fF
C1209 AdderSubtractor_0/XOR2IN_3/NAND2IN_1/w_n16_n4# AdderSubtractor_0/XOR2IN_3/NAND2IN_2/vin2 0.10fF
C1210 Enable_1/AND4Bit_1/AND2IN_2/NOT_0/in vdd 0.08fF
C1211 OR2IN_1/NOT_0/in gnd 0.11fF
C1212 AdderSubtractor_0/fullAdder_1/AND2IN_0/NOT_0/in AdderSubtractor_0/fullAdder_1/AND2IN_0/NAND2IN_0/w_n16_n4# 0.08fF
C1213 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_3/vin2 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_3/w_n16_n4# 0.10fF
C1214 Comparator_0/AND5IN_0/NOT_0/in vdd 0.37fF
C1215 AdderSubtractor_0/fullAdder_3/XOR2IN_1/vin1 AdderSubtractor_0/fullAdder_3/AND2IN_1/NOT_0/in 0.06fF
C1216 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_3/w_n16_n4# OR3IN_2/vin1 0.08fF
C1217 Enable_2/vinEn Enable_2/AND4Bit_1/AND2IN_2/NAND2IN_0/w_n16_n4# 0.10fF
C1218 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_0/w_n16_n4# AdderSubtractor_0/XOR2IN_1/vout 0.10fF
C1219 Decoder_0/AND4Bit_0/AND2IN_3/NOT_0/w_n7_n3# vdd 0.06fF
C1220 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_3/vin2 0.06fF
C1221 Comparator_0/XOR2IN_2/NAND2IN_2/vin2 vdd 0.08fF
C1222 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_1/w_n16_n4# vdd 0.11fF
C1223 AdderSubtractor_0/fullAdder_2/AND2IN_0/NOT_0/in AdderSubtractor_0/fullAdder_2/AND2IN_0/NAND2IN_0/w_n16_n4# 0.08fF
C1224 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_3/vin2 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_3/w_n16_n4# 0.10fF
C1225 OR3IN_1/NOT_0/in OR3IN_1/w_n19_n9# 0.05fF
C1226 Enable_2/AND4Bit_0/AND2IN_3/NOT_0/w_n7_n3# Enable_2/AND4Bit_0/AND2IN_3/NOT_0/in 0.07fF
C1227 Enable_1/AND4Bit_0/AND2IN_1/NAND2IN_0/w_n16_n4# vdd 0.11fF
C1228 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_3/w_n16_n4# AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_3/vin1 0.10fF
C1229 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_0/w_n16_n4# AdderSubtractor_0/XOR2IN_2/vout 0.10fF
C1230 vina1 vina2 3.01fF
C1231 AND4Bit_0/AND2IN_1/NOT_0/in Enable_2/voutb1 0.06fF
C1232 Comparator_0/AND2IN_1/NAND2IN_0/w_n16_n4# Comparator_0/AND4IN_0/vout 0.10fF
C1233 vdd AdderSubtractor_0/fullAdder_1/AND2IN_0/NAND2IN_0/w_n16_n4# 0.11fF
C1234 AdderSubtractor_0/XOR2IN_3/NAND2IN_2/vin2 AdderSubtractor_0/XOR2IN_3/NAND2IN_3/vin2 0.06fF
C1235 AdderSubtractor_0/fullAdder_2/AND2IN_0/NAND2IN_0/w_n16_n4# vdd 0.11fF
C1236 Comparator_0/XOR2IN_1/NAND2IN_1/w_n16_n4# vdd 0.11fF
C1237 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_1/w_n16_n4# AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_3/vin1 0.08fF
C1238 OR2IN_0/vout vina3 0.06fF
C1239 OR3IN_0/vin2 OR3IN_1/vin1 0.07fF
C1240 OR3IN_0/vin2 OR3IN_2/vin1 0.07fF
C1241 vdd AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_0/w_n16_n4# 0.11fF
C1242 vdd AdderSubtractor_0/fullAdder_1/AND2IN_1/NOT_0/w_n7_n3# 0.06fF
C1243 gnd AdderSubtractor_0/fullAdder_3/XOR2IN_1/vin1 0.52fF
C1244 Enable_1/vinEn Enable_1/AND4Bit_0/AND2IN_2/NAND2IN_0/w_n16_n4# 0.10fF
C1245 vina3 vinb3 0.19fF
C1246 AdderSubtractor_0/fullAdder_2/AND2IN_1/NOT_0/w_n7_n3# vdd 0.06fF
C1247 Comparator_0/XOR2IN_1/NAND2IN_3/vin2 vdd 0.08fF
C1248 Comparator_0/XOR2IN_0/NAND2IN_2/vin2 Comparator_0/XOR2IN_0/NAND2IN_3/vin2 0.06fF
C1249 Enable_2/AND4Bit_1/AND2IN_2/NOT_0/w_n7_n3# Enable_2/AND4Bit_1/AND2IN_2/NOT_0/in 0.07fF
C1250 OR2IN_0/vout vinb2 0.06fF
C1251 Comparator_0/NOT_5/out Comparator_0/NOT_4/out 0.14fF
C1252 Enable_1/voutb1 Comparator_0/NOT_2/w_n7_n3# 0.07fF
C1253 Comparator_0/NOT_0/out gnd 0.14fF
C1254 OR2IN_0/vin2 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_2/vin2 0.39fF
C1255 Enable_0/AND4Bit_0/AND2IN_1/NOT_0/w_n7_n3# Enable_0/vouta1 0.03fF
C1256 Comparator_0/NOT_2/out gnd 0.20fF
C1257 OR2IN_0/vin2 AdderSubtractor_0/XOR2IN_0/NAND2IN_2/vin2 0.39fF
C1258 Enable_2/AND4Bit_0/AND2IN_0/NOT_0/w_n7_n3# Enable_2/vouta0 0.03fF
C1259 Comparator_0/XOR2IN_3/NAND2IN_1/w_n16_n4# Comparator_0/XOR2IN_3/NAND2IN_2/vin2 0.10fF
C1260 Decoder_0/AND4Bit_0/AND2IN_0/NOT_0/w_n7_n3# OR2IN_0/vin1 0.03fF
C1261 Enable_2/vinEn Enable_2/AND4Bit_0/AND2IN_0/NOT_0/in 0.06fF
C1262 Enable_1/vouta0 Comparator_0/NOT_6/out 0.06fF
C1263 Comparator_0/AND2IN_1/NOT_0/w_n7_n3# OR3IN_0/vin2 0.03fF
C1264 Enable_2/AND4Bit_0/AND2IN_3/NOT_0/w_n7_n3# vdd 0.06fF
C1265 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_2/w_n16_n4# AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_3/vin2 0.08fF
C1266 vinb2 vinb3 1.72fF
C1267 Enable_1/voutb0 Comparator_0/NOT_3/w_n7_n3# 0.07fF
C1268 Enable_0/AND4Bit_0/AND2IN_3/NOT_0/w_n7_n3# Enable_0/vouta3 0.03fF
C1269 Comparator_0/XOR2IN_2/NAND2IN_3/vin1 gnd 0.13fF
C1270 AdderSubtractor_0/XOR2IN_0/NAND2IN_2/w_n16_n4# vdd 0.11fF
C1271 Comparator_0/NOT_5/out Enable_1/vouta3 0.06fF
C1272 Comparator_0/AND2IN_2/NAND2IN_0/w_n16_n4# Comparator_0/AND2IN_2/NOT_0/in 0.08fF
C1273 vdd Decoder_0/NOT_0/out 0.06fF
C1274 Enable_1/vouta3 Comparator_0/XOR2IN_3/NAND2IN_0/w_n16_n4# 0.10fF
C1275 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_0/w_n16_n4# 0.08fF
C1276 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_1/w_n16_n4# AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_3/vin1 0.08fF
C1277 Comparator_0/AND2IN_0/NOT_0/in gnd 0.05fF
C1278 AdderSubtractor_0/fullAdder_3/vcin AdderSubtractor_0/fullAdder_2/OR2IN_0/NOT_0/w_n7_n3# 0.03fF
C1279 AdderSubtractor_0/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/XOR2IN_1/NAND2IN_3/vin1 0.06fF
C1280 AdderSubtractor_0/fullAdder_2/vcin AdderSubtractor_0/fullAdder_2/XOR2IN_1/vin1 0.26fF
C1281 Enable_1/voutb3 gnd 0.29fF
C1282 Comparator_0/XOR2IN_3/NAND2IN_2/vin2 Comparator_0/XOR2IN_3/NAND2IN_3/vin2 0.06fF
C1283 Enable_2/AND4Bit_1/AND2IN_2/NOT_0/w_n7_n3# vdd 0.06fF
C1284 Enable_0/vouta2 AdderSubtractor_0/fullAdder_2/AND2IN_0/NAND2IN_0/w_n16_n4# 0.10fF
C1285 Enable_1/AND4Bit_0/AND2IN_3/NOT_0/w_n7_n3# Enable_1/AND4Bit_0/AND2IN_3/NOT_0/in 0.07fF
C1286 vdd Decoder_0/AND4Bit_0/AND2IN_0/NOT_0/in 0.08fF
C1287 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_3/vin2 OR3IN_2/vin1 0.06fF
C1288 Comparator_0/AND2IN_1/NOT_0/in vdd 0.08fF
C1289 Comparator_0/AND4IN_1/NOT_0/w_n7_n3# Comparator_0/AND4IN_1/NOT_0/in 0.07fF
C1290 Enable_2/AND4Bit_0/AND2IN_2/NAND2IN_0/w_n16_n4# vdd 0.11fF
C1291 AdderSubtractor_0/fullAdder_3/OR2IN_0/NOT_0/in AdderSubtractor_0/fullAdder_3/OR2IN_0/w_n19_n9# 0.05fF
C1292 vdd AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_2/w_n16_n4# 0.11fF
C1293 AdderSubtractor_0/XOR2IN_0/NAND2IN_3/vin1 vdd 0.43fF
C1294 OR2IN_0/w_n19_n9# vdd 0.09fF
C1295 vdd Decoder_0/AND4Bit_0/AND2IN_1/NOT_0/w_n7_n3# 0.06fF
C1296 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_2/w_n16_n4# vdd 0.11fF
C1297 gnd OR2IN_0/vin2 1.26fF
C1298 OR2IN_1/NOT_0/in OR2IN_1/vin2 0.08fF
C1299 OR2IN_1/NOT_0/w_n7_n3# vdd 0.06fF
C1300 gnd AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_2/vin2 0.19fF
C1301 gnd AdderSubtractor_0/XOR2IN_0/NAND2IN_2/vin2 0.19fF
C1302 gnd AdderSubtractor_0/fullAdder_3/AND2IN_1/NOT_0/in 0.05fF
C1303 Enable_0/voutb2 Enable_0/voutb3 3.36fF
C1304 OR2IN_0/vout Enable_0/AND4Bit_1/AND2IN_0/NAND2IN_0/w_n16_n4# 0.10fF
C1305 AND4Bit_0/AND2IN_0/NAND2IN_0/w_n16_n4# AND4Bit_0/AND2IN_0/NOT_0/in 0.08fF
C1306 Enable_1/voutb2 Comparator_0/XOR2IN_2/NAND2IN_2/w_n16_n4# 0.10fF
C1307 OR3IN_0/w_n19_n9# OR3IN_0/NOT_0/in 0.05fF
C1308 AdderSubtractor_0/XOR2IN_1/NAND2IN_0/w_n16_n4# AdderSubtractor_0/XOR2IN_1/NAND2IN_2/vin2 0.08fF
C1309 vina2 Enable_2/vinEn 0.19fF
C1310 Comparator_0/NOT_6/out Comparator_0/NOT_3/out 0.06fF
C1311 Enable_1/vinEn Enable_1/AND4Bit_0/AND2IN_0/NAND2IN_0/w_n16_n4# 0.10fF
C1312 vdd AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_2/w_n16_n4# 0.11fF
C1313 Enable_1/AND4Bit_1/AND2IN_2/NOT_0/w_n7_n3# Enable_1/AND4Bit_1/AND2IN_2/NOT_0/in 0.07fF
C1314 AND4Bit_0/AND2IN_1/NOT_0/in AND4Bit_0/AND2IN_1/NAND2IN_0/w_n16_n4# 0.08fF
C1315 Comparator_0/AND5IN_0/w_n26_1# Comparator_0/NOT_6/out 0.12fF
C1316 gnd Enable_2/AND4Bit_1/AND2IN_3/NOT_0/in 0.05fF
C1317 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_3/w_n16_n4# vdd 0.11fF
C1318 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_2/w_n16_n4# AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_2/vin2 0.10fF
C1319 Enable_0/AND4Bit_0/AND2IN_3/NOT_0/w_n7_n3# vdd 0.06fF
C1320 Comparator_0/XOR2IN_3/NAND2IN_3/vin1 vdd 0.43fF
C1321 Comparator_0/XOR2IN_1/NAND2IN_2/vin2 Comparator_0/XOR2IN_1/NAND2IN_3/vin1 0.06fF
C1322 vout2 OR3IN_1/vin3 0.06fF
C1323 Enable_1/vinEn Enable_1/AND4Bit_1/AND2IN_3/NAND2IN_0/w_n16_n4# 0.10fF
C1324 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_3/w_n16_n4# AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_3/vin1 0.10fF
C1325 vina0 gnd 0.19fF
C1326 OR3IN_0/vin3 OR3IN_0/vin2 0.14fF
C1327 Decoder_0/AND4Bit_0/AND2IN_2/NAND2IN_0/w_n16_n4# vinSel1 0.10fF
C1328 OR3IN_2/vin3 vdd 0.25fF
C1329 vdd AdderSubtractor_0/fullAdder_1/OR2IN_0/NOT_0/w_n7_n3# 0.06fF
C1330 OR2IN_0/vin2 AdderSubtractor_0/XOR2IN_1/vout 0.06fF
C1331 OR2IN_0/vin2 AdderSubtractor_0/XOR2IN_3/NAND2IN_2/vin2 0.39fF
C1332 AdderSubtractor_0/fullAdder_2/OR2IN_0/NOT_0/w_n7_n3# vdd 0.06fF
C1333 Enable_0/AND4Bit_1/AND2IN_2/NOT_0/w_n7_n3# vdd 0.06fF
C1334 AdderSubtractor_0/XOR2IN_2/vout OR2IN_0/vin2 0.06fF
C1335 AdderSubtractor_0/fullAdder_3/vcin AdderSubtractor_0/XOR2IN_3/vout 0.06fF
C1336 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_3/vin2 OR2IN_1/vin1 0.06fF
C1337 Enable_1/AND4Bit_1/AND2IN_1/NAND2IN_0/w_n16_n4# vdd 0.11fF
C1338 gnd AdderSubtractor_0/fullAdder_3/AND2IN_0/NOT_0/in 0.05fF
C1339 Enable_0/AND4Bit_0/AND2IN_3/NOT_0/w_n7_n3# Enable_0/AND4Bit_0/AND2IN_3/NOT_0/in 0.07fF
C1340 OR3IN_0/w_n19_n9# vdd 0.10fF
C1341 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_2/vin2 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_2/w_n16_n4# 0.10fF
C1342 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_1/w_n16_n4# vdd 0.11fF
C1343 Comparator_0/AND3IN_0/NOT_0/in vdd 0.19fF
C1344 Enable_0/vouta3 AdderSubtractor_0/XOR2IN_3/vout 0.27fF
C1345 Enable_2/AND4Bit_0/AND2IN_0/NAND2IN_0/w_n16_n4# vdd 0.11fF
C1346 AND4Bit_0/AND2IN_1/NOT_0/w_n7_n3# AND4Bit_0/AND2IN_1/NOT_0/in 0.07fF
C1347 AND4Bit_0/AND2IN_3/NOT_0/w_n7_n3# OR2IN_1/vin2 0.03fF
C1348 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_2/w_n16_n4# AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_2/vin2 0.10fF
C1349 Comparator_0/NOT_5/out vdd 0.12fF
C1350 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_2/vin2 vdd 0.15fF
C1351 Comparator_0/XOR2IN_3/NAND2IN_0/w_n16_n4# vdd 0.11fF
C1352 Comparator_0/XOR2IN_1/NAND2IN_0/w_n16_n4# Comparator_0/XOR2IN_1/NAND2IN_2/vin2 0.08fF
C1353 AdderSubtractor_0/fullAdder_2/XOR2IN_1/vin1 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_3/w_n16_n4# 0.08fF
C1354 Comparator_0/OR4IN_0/vin1 vdd 0.21fF
C1355 OR2IN_0/vout Enable_0/AND4Bit_1/AND2IN_0/NOT_0/in 0.06fF
C1356 gnd AdderSubtractor_0/fullAdder_1/OR2IN_0/vin1 0.26fF
C1357 Decoder_0/AND4Bit_0/AND2IN_3/NOT_0/in vdd 0.08fF
C1358 gnd AdderSubtractor_0/fullAdder_3/OR2IN_0/vin2 0.27fF
C1359 Decoder_0/AND4Bit_0/AND2IN_2/NOT_0/in Decoder_0/AND4Bit_0/AND2IN_2/NOT_0/w_n7_n3# 0.07fF
C1360 gnd AdderSubtractor_0/fullAdder_2/OR2IN_0/vin1 0.26fF
C1361 Enable_2/AND4Bit_1/AND2IN_3/NAND2IN_0/w_n16_n4# vdd 0.11fF
C1362 gnd AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_3/vin1 0.06fF
C1363 OR3IN_1/w_n19_n9# vdd 0.10fF
C1364 gnd AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_3/vin1 0.06fF
C1365 OR3IN_0/vin2 OR3IN_1/vin2 4.88fF
C1366 vina1 Enable_2/AND4Bit_0/AND2IN_1/NAND2IN_0/w_n16_n4# 0.10fF
C1367 Enable_0/AND4Bit_1/AND2IN_2/NOT_0/w_n7_n3# Enable_0/AND4Bit_1/AND2IN_2/NOT_0/in 0.07fF
C1368 gnd Enable_0/AND4Bit_1/AND2IN_3/NOT_0/in 0.05fF
C1369 Enable_1/vouta1 Comparator_0/NOT_6/out 0.06fF
C1370 gnd AdderSubtractor_0/XOR2IN_1/vout 0.28fF
C1371 AdderSubtractor_0/fullAdder_0/XOR2IN_1/vin1 AdderSubtractor_0/fullAdder_0/AND2IN_1/NAND2IN_0/w_n16_n4# 0.10fF
C1372 AdderSubtractor_0/XOR2IN_0/vout AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_2/vin2 0.39fF
C1373 Enable_1/vinEn vinb3 0.13fF
C1374 gnd AdderSubtractor_0/XOR2IN_3/NAND2IN_2/vin2 0.19fF
C1375 gnd Enable_2/vouta3 0.14fF
C1376 gnd AdderSubtractor_0/XOR2IN_2/vout 0.28fF
C1377 Comparator_0/AND3IN_0/NOT_0/w_n7_n3# Comparator_0/OR4IN_0/vin2 0.03fF
C1378 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_3/vin2 vdd 0.08fF
C1379 OR3IN_0/vin2 OR3IN_2/vin2 0.11fF
C1380 gnd Decoder_0/AND4Bit_0/AND2IN_1/NOT_0/in 0.05fF
C1381 AdderSubtractor_0/XOR2IN_0/NAND2IN_3/vin2 vdd 0.08fF
C1382 AdderSubtractor_0/XOR2IN_2/vout AdderSubtractor_0/XOR2IN_2/NAND2IN_3/w_n16_n4# 0.08fF
C1383 AdderSubtractor_0/fullAdder_3/OR2IN_0/vin1 vdd 0.06fF
C1384 Enable_1/voutb3 Enable_1/AND4Bit_1/AND2IN_3/NOT_0/w_n7_n3# 0.03fF
C1385 gnd AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_2/vin2 0.19fF
C1386 Enable_1/vouta0 Enable_1/vinEn 23.23fF
C1387 Comparator_0/XOR2IN_0/NAND2IN_2/vin2 gnd 0.19fF
C1388 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_3/vin1 vdd 0.43fF
C1389 gnd Enable_2/voutb2 0.14fF
C1390 AdderSubtractor_0/XOR2IN_3/NAND2IN_3/w_n16_n4# vdd 0.11fF
C1391 AdderSubtractor_0/fullAdder_3/OR2IN_0/w_n19_n9# vdd 0.09fF
C1392 Enable_1/vinEn Comparator_0/AND2IN_2/NAND2IN_0/w_n16_n4# 0.10fF
C1393 AdderSubtractor_0/fullAdder_1/OR2IN_0/vin1 AdderSubtractor_0/fullAdder_1/OR2IN_0/w_n19_n9# 0.16fF
C1394 AdderSubtractor_0/XOR2IN_3/vout vdd 0.20fF
C1395 AdderSubtractor_0/fullAdder_3/XOR2IN_1/vin1 AdderSubtractor_0/fullAdder_3/AND2IN_1/NAND2IN_0/w_n16_n4# 0.10fF
C1396 gnd AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_3/vin1 0.06fF
C1397 Enable_2/voutb3 vdd 0.06fF
C1398 gnd Enable_2/AND4Bit_0/AND2IN_0/NOT_0/in 0.05fF
C1399 Enable_1/AND4Bit_0/AND2IN_0/NOT_0/w_n7_n3# vdd 0.06fF
C1400 Comparator_0/NOT_5/out Comparator_0/NOT_4/in 0.06fF
C1401 vout3 gnd 0.07fF
C1402 AND4Bit_0/AND2IN_0/NAND2IN_0/w_n16_n4# vdd 0.11fF
C1403 AdderSubtractor_0/XOR2IN_0/NAND2IN_3/vin2 AdderSubtractor_0/XOR2IN_0/vout 0.06fF
C1404 gnd AdderSubtractor_0/XOR2IN_2/NAND2IN_3/vin2 0.06fF
C1405 AdderSubtractor_0/fullAdder_2/OR2IN_0/vin1 AdderSubtractor_0/fullAdder_2/OR2IN_0/w_n19_n9# 0.16fF
C1406 Comparator_0/XOR2IN_0/NAND2IN_3/w_n16_n4# vdd 0.11fF
C1407 Comparator_0/XOR2IN_0/NAND2IN_0/w_n16_n4# Enable_1/vouta0 0.10fF
C1408 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_2/vin2 vdd 0.08fF
C1409 Comparator_0/NOT_3/w_n7_n3# vdd 0.06fF
C1410 Enable_0/voutb2 OR2IN_0/vin2 0.06fF
C1411 Comparator_0/XOR2IN_2/NAND2IN_2/w_n16_n4# vdd 0.11fF
C1412 Enable_0/vouta0 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_1/w_n16_n4# 0.10fF
C1413 gnd OR2IN_1/vin2 0.19fF
C1414 AdderSubtractor_0/XOR2IN_2/NAND2IN_3/vin2 AdderSubtractor_0/XOR2IN_2/NAND2IN_3/w_n16_n4# 0.10fF
C1415 OR2IN_0/NOT_0/in OR2IN_0/w_n19_n9# 0.05fF
C1416 AdderSubtractor_0/XOR2IN_3/NAND2IN_2/w_n16_n4# AdderSubtractor_0/XOR2IN_3/NAND2IN_3/vin2 0.08fF
C1417 Decoder_0/AND4Bit_0/AND2IN_2/NOT_0/in gnd 0.05fF
C1418 vdd AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_3/vin1 0.43fF
C1419 Enable_0/AND4Bit_1/AND2IN_3/NAND2IN_0/w_n16_n4# vdd 0.11fF
C1420 AdderSubtractor_0/fullAdder_2/XOR2IN_1/vin1 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_3/vin2 0.06fF
C1421 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_3/vin1 vdd 0.43fF
C1422 Enable_1/voutb2 Comparator_0/NOT_2/out 0.06fF
C1423 Comparator_0/NOR2IN_0/w_n19_n9# OR3IN_2/vin2 0.12fF
C1424 Decoder_0/NOT_1/out Decoder_0/NOT_0/out 0.99fF
C1425 vina3 vinb1 0.19fF
C1426 Enable_0/vouta1 AdderSubtractor_0/fullAdder_1/AND2IN_0/NAND2IN_0/w_n16_n4# 0.10fF
C1427 Enable_2/vinEn Enable_2/AND4Bit_0/AND2IN_3/NOT_0/in 0.06fF
C1428 Enable_1/vinEn Comparator_0/AND4IN_0/vout 0.06fF
C1429 Comparator_0/AND3IN_0/NOT_0/in Comparator_0/NOT_1/out 0.06fF
C1430 OR3IN_0/vin3 vcout 0.06fF
C1431 AdderSubtractor_0/fullAdder_1/vcin AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_0/w_n16_n4# 0.10fF
C1432 Enable_1/vinEn OR3IN_2/vin2 0.06fF
C1433 Comparator_0/NOT_0/out Comparator_0/NOT_4/out 0.06fF
C1434 Enable_2/vouta3 Enable_2/voutb2 0.06fF
C1435 gnd AdderSubtractor_0/fullAdder_2/OR2IN_0/vin2 0.27fF
C1436 Comparator_0/NOT_2/out Comparator_0/NOT_4/out 0.06fF
C1437 Comparator_0/NOT_5/in gnd 0.07fF
C1438 Comparator_0/NOT_5/out Comparator_0/NOT_1/out 0.06fF
C1439 vinb1 vinb2 1.72fF
C1440 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_3/vin2 vdd 0.08fF
C1441 Comparator_0/XOR2IN_1/NAND2IN_2/vin2 vdd 0.08fF
C1442 AdderSubtractor_0/XOR2IN_3/NAND2IN_1/w_n16_n4# vdd 0.11fF
C1443 Enable_2/vinEn Enable_2/AND4Bit_1/AND2IN_2/NOT_0/in 0.06fF
C1444 Enable_1/voutb2 Enable_1/voutb3 15.34fF
C1445 Comparator_0/XOR2IN_0/NAND2IN_2/w_n16_n4# Comparator_0/XOR2IN_0/NAND2IN_3/vin2 0.08fF
C1446 vina0 vina2 0.19fF
C1447 AdderSubtractor_0/fullAdder_1/OR2IN_0/w_n19_n9# Gnd 1.40fF
C1448 AdderSubtractor_0/fullAdder_1/OR2IN_0/NOT_0/in Gnd 0.42fF
C1449 AdderSubtractor_0/fullAdder_1/OR2IN_0/NOT_0/w_n7_n3# Gnd 0.61fF
C1450 AdderSubtractor_0/fullAdder_1/AND2IN_1/NOT_0/in Gnd 0.37fF
C1451 AdderSubtractor_0/fullAdder_1/AND2IN_1/NOT_0/w_n7_n3# Gnd 0.61fF
C1452 AdderSubtractor_0/fullAdder_1/XOR2IN_1/vin1 Gnd 3.73fF
C1453 AdderSubtractor_0/fullAdder_1/AND2IN_1/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1454 AdderSubtractor_0/fullAdder_1/AND2IN_0/NOT_0/in Gnd 0.37fF
C1455 AdderSubtractor_0/fullAdder_1/AND2IN_0/NOT_0/w_n7_n3# Gnd 0.61fF
C1456 AdderSubtractor_0/fullAdder_1/AND2IN_0/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1457 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_3/vin1 Gnd 0.54fF
C1458 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_3/w_n16_n4# Gnd 1.16fF
C1459 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_3/vin2 Gnd 0.55fF
C1460 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_2/vin2 Gnd 0.80fF
C1461 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_2/w_n16_n4# Gnd 1.16fF
C1462 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_1/w_n16_n4# Gnd 1.16fF
C1463 AdderSubtractor_0/XOR2IN_1/vout Gnd 6.27fF
C1464 Enable_0/vouta1 Gnd 15.71fF
C1465 AdderSubtractor_0/fullAdder_1/XOR2IN_0/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1466 OR3IN_1/vin1 Gnd 2.25fF
C1467 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_3/vin1 Gnd 0.54fF
C1468 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_3/w_n16_n4# Gnd 1.16fF
C1469 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_3/vin2 Gnd 0.55fF
C1470 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_2/vin2 Gnd 0.80fF
C1471 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_2/w_n16_n4# Gnd 1.16fF
C1472 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_1/w_n16_n4# Gnd 1.16fF
C1473 AdderSubtractor_0/fullAdder_1/vcin Gnd 6.72fF
C1474 AdderSubtractor_0/fullAdder_1/XOR2IN_1/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1475 AdderSubtractor_0/fullAdder_0/OR2IN_0/w_n19_n9# Gnd 1.40fF
C1476 AdderSubtractor_0/fullAdder_0/OR2IN_0/NOT_0/in Gnd 0.42fF
C1477 AdderSubtractor_0/fullAdder_0/OR2IN_0/NOT_0/w_n7_n3# Gnd 0.61fF
C1478 AdderSubtractor_0/fullAdder_0/AND2IN_1/NOT_0/in Gnd 0.37fF
C1479 AdderSubtractor_0/fullAdder_0/AND2IN_1/NOT_0/w_n7_n3# Gnd 0.61fF
C1480 AdderSubtractor_0/fullAdder_0/XOR2IN_1/vin1 Gnd 3.73fF
C1481 AdderSubtractor_0/fullAdder_0/AND2IN_1/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1482 vdd Gnd 38.37fF
C1483 AdderSubtractor_0/fullAdder_0/AND2IN_0/NOT_0/in Gnd 0.37fF
C1484 AdderSubtractor_0/fullAdder_0/AND2IN_0/NOT_0/w_n7_n3# Gnd 0.61fF
C1485 AdderSubtractor_0/fullAdder_0/AND2IN_0/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1486 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_3/vin1 Gnd 0.54fF
C1487 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_3/w_n16_n4# Gnd 1.16fF
C1488 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_3/vin2 Gnd 0.55fF
C1489 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_2/vin2 Gnd 0.80fF
C1490 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_2/w_n16_n4# Gnd 1.16fF
C1491 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_1/w_n16_n4# Gnd 1.16fF
C1492 AdderSubtractor_0/XOR2IN_0/vout Gnd 3.62fF
C1493 Enable_0/vouta0 Gnd 9.74fF
C1494 AdderSubtractor_0/fullAdder_0/XOR2IN_0/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1495 OR3IN_0/vin1 Gnd 1.16fF
C1496 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_3/vin1 Gnd 0.54fF
C1497 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_3/w_n16_n4# Gnd 1.16fF
C1498 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_3/vin2 Gnd 0.55fF
C1499 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_2/vin2 Gnd 0.80fF
C1500 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_2/w_n16_n4# Gnd 1.16fF
C1501 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_1/w_n16_n4# Gnd 1.16fF
C1502 AdderSubtractor_0/fullAdder_0/XOR2IN_1/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1503 AdderSubtractor_0/XOR2IN_3/NAND2IN_3/vin1 Gnd 0.54fF
C1504 AdderSubtractor_0/XOR2IN_3/NAND2IN_3/w_n16_n4# Gnd 1.16fF
C1505 AdderSubtractor_0/XOR2IN_3/NAND2IN_3/vin2 Gnd 0.55fF
C1506 AdderSubtractor_0/XOR2IN_3/NAND2IN_2/vin2 Gnd 0.80fF
C1507 AdderSubtractor_0/XOR2IN_3/NAND2IN_2/w_n16_n4# Gnd 1.16fF
C1508 AdderSubtractor_0/XOR2IN_3/NAND2IN_1/w_n16_n4# Gnd 1.16fF
C1509 AdderSubtractor_0/XOR2IN_3/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1510 AdderSubtractor_0/XOR2IN_2/NAND2IN_3/vin1 Gnd 0.54fF
C1511 AdderSubtractor_0/XOR2IN_2/NAND2IN_3/w_n16_n4# Gnd 1.16fF
C1512 AdderSubtractor_0/XOR2IN_2/NAND2IN_3/vin2 Gnd 0.55fF
C1513 AdderSubtractor_0/XOR2IN_2/NAND2IN_2/vin2 Gnd 0.80fF
C1514 AdderSubtractor_0/XOR2IN_2/NAND2IN_2/w_n16_n4# Gnd 1.16fF
C1515 AdderSubtractor_0/XOR2IN_2/NAND2IN_1/w_n16_n4# Gnd 1.16fF
C1516 AdderSubtractor_0/XOR2IN_2/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1517 AdderSubtractor_0/XOR2IN_1/NAND2IN_3/vin1 Gnd 0.54fF
C1518 AdderSubtractor_0/XOR2IN_1/NAND2IN_3/w_n16_n4# Gnd 1.16fF
C1519 AdderSubtractor_0/XOR2IN_1/NAND2IN_3/vin2 Gnd 0.55fF
C1520 AdderSubtractor_0/XOR2IN_1/NAND2IN_2/vin2 Gnd 0.80fF
C1521 AdderSubtractor_0/XOR2IN_1/NAND2IN_2/w_n16_n4# Gnd 1.16fF
C1522 AdderSubtractor_0/XOR2IN_1/NAND2IN_1/w_n16_n4# Gnd 1.16fF
C1523 AdderSubtractor_0/XOR2IN_1/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1524 AdderSubtractor_0/XOR2IN_0/NAND2IN_3/vin1 Gnd 0.54fF
C1525 AdderSubtractor_0/XOR2IN_0/NAND2IN_3/w_n16_n4# Gnd 1.16fF
C1526 AdderSubtractor_0/XOR2IN_0/NAND2IN_3/vin2 Gnd 0.55fF
C1527 AdderSubtractor_0/XOR2IN_0/NAND2IN_2/vin2 Gnd 0.80fF
C1528 AdderSubtractor_0/XOR2IN_0/NAND2IN_2/w_n16_n4# Gnd 1.16fF
C1529 AdderSubtractor_0/XOR2IN_0/NAND2IN_1/w_n16_n4# Gnd 1.16fF
C1530 OR2IN_0/vin2 Gnd 21.96fF
C1531 AdderSubtractor_0/XOR2IN_0/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1532 AdderSubtractor_0/fullAdder_3/OR2IN_0/w_n19_n9# Gnd 1.40fF
C1533 vcout Gnd 0.22fF
C1534 AdderSubtractor_0/fullAdder_3/OR2IN_0/NOT_0/in Gnd 0.42fF
C1535 AdderSubtractor_0/fullAdder_3/OR2IN_0/NOT_0/w_n7_n3# Gnd 0.61fF
C1536 AdderSubtractor_0/fullAdder_3/AND2IN_1/NOT_0/in Gnd 0.37fF
C1537 AdderSubtractor_0/fullAdder_3/AND2IN_1/NOT_0/w_n7_n3# Gnd 0.61fF
C1538 AdderSubtractor_0/fullAdder_3/XOR2IN_1/vin1 Gnd 3.73fF
C1539 AdderSubtractor_0/fullAdder_3/AND2IN_1/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1540 AdderSubtractor_0/fullAdder_3/AND2IN_0/NOT_0/in Gnd 0.37fF
C1541 AdderSubtractor_0/fullAdder_3/AND2IN_0/NOT_0/w_n7_n3# Gnd 0.61fF
C1542 AdderSubtractor_0/fullAdder_3/AND2IN_0/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1543 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_3/vin1 Gnd 0.54fF
C1544 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_3/w_n16_n4# Gnd 1.16fF
C1545 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_3/vin2 Gnd 0.55fF
C1546 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_2/vin2 Gnd 0.80fF
C1547 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_2/w_n16_n4# Gnd 1.16fF
C1548 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_1/w_n16_n4# Gnd 1.16fF
C1549 AdderSubtractor_0/XOR2IN_3/vout Gnd 6.38fF
C1550 Enable_0/vouta3 Gnd 20.73fF
C1551 AdderSubtractor_0/fullAdder_3/XOR2IN_0/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1552 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_3/vin1 Gnd 0.54fF
C1553 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_3/w_n16_n4# Gnd 1.16fF
C1554 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_3/vin2 Gnd 0.55fF
C1555 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_2/vin2 Gnd 0.80fF
C1556 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_2/w_n16_n4# Gnd 1.16fF
C1557 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_1/w_n16_n4# Gnd 1.16fF
C1558 AdderSubtractor_0/fullAdder_3/vcin Gnd 6.69fF
C1559 AdderSubtractor_0/fullAdder_3/XOR2IN_1/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1560 AdderSubtractor_0/fullAdder_2/OR2IN_0/w_n19_n9# Gnd 1.40fF
C1561 AdderSubtractor_0/fullAdder_2/OR2IN_0/NOT_0/in Gnd 0.42fF
C1562 AdderSubtractor_0/fullAdder_2/OR2IN_0/NOT_0/w_n7_n3# Gnd 0.61fF
C1563 AdderSubtractor_0/fullAdder_2/AND2IN_1/NOT_0/in Gnd 0.37fF
C1564 AdderSubtractor_0/fullAdder_2/AND2IN_1/NOT_0/w_n7_n3# Gnd 0.61fF
C1565 AdderSubtractor_0/fullAdder_2/XOR2IN_1/vin1 Gnd 3.73fF
C1566 AdderSubtractor_0/fullAdder_2/AND2IN_1/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1567 AdderSubtractor_0/fullAdder_2/AND2IN_0/NOT_0/in Gnd 0.37fF
C1568 AdderSubtractor_0/fullAdder_2/AND2IN_0/NOT_0/w_n7_n3# Gnd 0.61fF
C1569 AdderSubtractor_0/fullAdder_2/AND2IN_0/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1570 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_3/vin1 Gnd 0.54fF
C1571 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_3/w_n16_n4# Gnd 1.16fF
C1572 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_3/vin2 Gnd 0.55fF
C1573 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_2/vin2 Gnd 0.80fF
C1574 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_2/w_n16_n4# Gnd 1.16fF
C1575 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_1/w_n16_n4# Gnd 1.16fF
C1576 AdderSubtractor_0/XOR2IN_2/vout Gnd 6.48fF
C1577 Enable_0/vouta2 Gnd 18.42fF
C1578 AdderSubtractor_0/fullAdder_2/XOR2IN_0/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1579 OR3IN_2/vin1 Gnd 1.40fF
C1580 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_3/vin1 Gnd 0.54fF
C1581 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_3/w_n16_n4# Gnd 1.16fF
C1582 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_3/vin2 Gnd 0.55fF
C1583 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_2/vin2 Gnd 0.80fF
C1584 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_2/w_n16_n4# Gnd 1.16fF
C1585 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_1/w_n16_n4# Gnd 1.16fF
C1586 AdderSubtractor_0/fullAdder_2/vcin Gnd 6.68fF
C1587 AdderSubtractor_0/fullAdder_2/XOR2IN_1/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1588 Enable_2/AND4Bit_1/AND2IN_3/NOT_0/in Gnd 0.37fF
C1589 Enable_2/AND4Bit_1/AND2IN_3/NOT_0/w_n7_n3# Gnd 0.61fF
C1590 Enable_2/AND4Bit_1/AND2IN_3/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1591 Enable_2/voutb2 Gnd 0.93fF
C1592 Enable_2/AND4Bit_1/AND2IN_2/NOT_0/in Gnd 0.37fF
C1593 Enable_2/AND4Bit_1/AND2IN_2/NOT_0/w_n7_n3# Gnd 0.61fF
C1594 Enable_2/AND4Bit_1/AND2IN_2/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1595 Enable_2/AND4Bit_1/AND2IN_1/NOT_0/in Gnd 0.37fF
C1596 Enable_2/AND4Bit_1/AND2IN_1/NOT_0/w_n7_n3# Gnd 0.61fF
C1597 Enable_2/AND4Bit_1/AND2IN_1/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1598 Enable_2/AND4Bit_1/AND2IN_0/NOT_0/in Gnd 0.37fF
C1599 Enable_2/AND4Bit_1/AND2IN_0/NOT_0/w_n7_n3# Gnd 0.61fF
C1600 Enable_2/AND4Bit_1/AND2IN_0/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1601 Enable_2/vouta3 Gnd 0.66fF
C1602 Enable_2/AND4Bit_0/AND2IN_3/NOT_0/in Gnd 0.37fF
C1603 Enable_2/AND4Bit_0/AND2IN_3/NOT_0/w_n7_n3# Gnd 0.61fF
C1604 Enable_2/AND4Bit_0/AND2IN_3/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1605 Enable_2/AND4Bit_0/AND2IN_2/NOT_0/in Gnd 0.37fF
C1606 Enable_2/AND4Bit_0/AND2IN_2/NOT_0/w_n7_n3# Gnd 0.61fF
C1607 Enable_2/AND4Bit_0/AND2IN_2/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1608 Enable_2/AND4Bit_0/AND2IN_1/NOT_0/in Gnd 0.37fF
C1609 Enable_2/AND4Bit_0/AND2IN_1/NOT_0/w_n7_n3# Gnd 0.61fF
C1610 Enable_2/AND4Bit_0/AND2IN_1/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1611 Enable_2/AND4Bit_0/AND2IN_0/NOT_0/in Gnd 0.37fF
C1612 Enable_2/AND4Bit_0/AND2IN_0/NOT_0/w_n7_n3# Gnd 0.61fF
C1613 Enable_2/vinEn Gnd 3.76fF
C1614 Enable_2/AND4Bit_0/AND2IN_0/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1615 Enable_1/AND4Bit_1/AND2IN_3/NOT_0/in Gnd 0.37fF
C1616 Enable_1/AND4Bit_1/AND2IN_3/NOT_0/w_n7_n3# Gnd 0.61fF
C1617 Enable_1/AND4Bit_1/AND2IN_3/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1618 Enable_1/AND4Bit_1/AND2IN_2/NOT_0/in Gnd 0.37fF
C1619 Enable_1/AND4Bit_1/AND2IN_2/NOT_0/w_n7_n3# Gnd 0.61fF
C1620 Enable_1/AND4Bit_1/AND2IN_2/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1621 Enable_1/AND4Bit_1/AND2IN_1/NOT_0/in Gnd 0.37fF
C1622 Enable_1/AND4Bit_1/AND2IN_1/NOT_0/w_n7_n3# Gnd 0.61fF
C1623 Enable_1/AND4Bit_1/AND2IN_1/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1624 Enable_1/AND4Bit_1/AND2IN_0/NOT_0/in Gnd 0.37fF
C1625 Enable_1/AND4Bit_1/AND2IN_0/NOT_0/w_n7_n3# Gnd 0.61fF
C1626 Enable_1/AND4Bit_1/AND2IN_0/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1627 Enable_1/AND4Bit_0/AND2IN_3/NOT_0/in Gnd 0.37fF
C1628 Enable_1/AND4Bit_0/AND2IN_3/NOT_0/w_n7_n3# Gnd 0.61fF
C1629 Enable_1/AND4Bit_0/AND2IN_3/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1630 Enable_1/AND4Bit_0/AND2IN_2/NOT_0/in Gnd 0.37fF
C1631 Enable_1/AND4Bit_0/AND2IN_2/NOT_0/w_n7_n3# Gnd 0.61fF
C1632 Enable_1/AND4Bit_0/AND2IN_2/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1633 Enable_1/AND4Bit_0/AND2IN_1/NOT_0/in Gnd 0.37fF
C1634 Enable_1/AND4Bit_0/AND2IN_1/NOT_0/w_n7_n3# Gnd 0.61fF
C1635 Enable_1/AND4Bit_0/AND2IN_1/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1636 Enable_1/AND4Bit_0/AND2IN_0/NOT_0/in Gnd 0.37fF
C1637 Enable_1/AND4Bit_0/AND2IN_0/NOT_0/w_n7_n3# Gnd 0.61fF
C1638 Enable_1/vinEn Gnd 30.92fF
C1639 Enable_1/AND4Bit_0/AND2IN_0/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1640 Enable_0/voutb3 Gnd 12.54fF
C1641 Enable_0/AND4Bit_1/AND2IN_3/NOT_0/in Gnd 0.37fF
C1642 Enable_0/AND4Bit_1/AND2IN_3/NOT_0/w_n7_n3# Gnd 0.61fF
C1643 vinb3 Gnd 23.79fF
C1644 Enable_0/AND4Bit_1/AND2IN_3/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1645 Enable_0/voutb2 Gnd 22.27fF
C1646 Enable_0/AND4Bit_1/AND2IN_2/NOT_0/in Gnd 0.37fF
C1647 Enable_0/AND4Bit_1/AND2IN_2/NOT_0/w_n7_n3# Gnd 0.61fF
C1648 vinb2 Gnd 23.90fF
C1649 Enable_0/AND4Bit_1/AND2IN_2/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1650 Enable_0/voutb1 Gnd 13.25fF
C1651 Enable_0/AND4Bit_1/AND2IN_1/NOT_0/in Gnd 0.37fF
C1652 Enable_0/AND4Bit_1/AND2IN_1/NOT_0/w_n7_n3# Gnd 0.61fF
C1653 vinb1 Gnd 24.00fF
C1654 Enable_0/AND4Bit_1/AND2IN_1/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1655 Enable_0/voutb0 Gnd 0.08fF
C1656 Enable_0/AND4Bit_1/AND2IN_0/NOT_0/in Gnd 0.37fF
C1657 Enable_0/AND4Bit_1/AND2IN_0/NOT_0/w_n7_n3# Gnd 0.61fF
C1658 vinb0 Gnd 24.10fF
C1659 Enable_0/AND4Bit_1/AND2IN_0/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1660 Enable_0/AND4Bit_0/AND2IN_3/NOT_0/in Gnd 0.37fF
C1661 Enable_0/AND4Bit_0/AND2IN_3/NOT_0/w_n7_n3# Gnd 0.61fF
C1662 vina3 Gnd 24.19fF
C1663 Enable_0/AND4Bit_0/AND2IN_3/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1664 Enable_0/AND4Bit_0/AND2IN_2/NOT_0/in Gnd 0.37fF
C1665 Enable_0/AND4Bit_0/AND2IN_2/NOT_0/w_n7_n3# Gnd 0.61fF
C1666 vina2 Gnd 24.29fF
C1667 Enable_0/AND4Bit_0/AND2IN_2/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1668 Enable_0/AND4Bit_0/AND2IN_1/NOT_0/in Gnd 0.37fF
C1669 Enable_0/AND4Bit_0/AND2IN_1/NOT_0/w_n7_n3# Gnd 0.61fF
C1670 vina1 Gnd 24.38fF
C1671 Enable_0/AND4Bit_0/AND2IN_1/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1672 gnd Gnd 42.07fF
C1673 Enable_0/AND4Bit_0/AND2IN_0/NOT_0/in Gnd 0.37fF
C1674 Enable_0/AND4Bit_0/AND2IN_0/NOT_0/w_n7_n3# Gnd 0.61fF
C1675 OR2IN_0/vout Gnd 3.38fF
C1676 vina0 Gnd 24.44fF
C1677 Enable_0/AND4Bit_0/AND2IN_0/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1678 OR2IN_1/vin2 Gnd 1.00fF
C1679 AND4Bit_0/AND2IN_3/NOT_0/in Gnd 0.37fF
C1680 AND4Bit_0/AND2IN_3/NOT_0/w_n7_n3# Gnd 0.61fF
C1681 AND4Bit_0/AND2IN_3/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1682 OR3IN_2/vin3 Gnd 1.28fF
C1683 AND4Bit_0/AND2IN_2/NOT_0/in Gnd 0.37fF
C1684 AND4Bit_0/AND2IN_2/NOT_0/w_n7_n3# Gnd 0.61fF
C1685 AND4Bit_0/AND2IN_2/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1686 OR3IN_1/vin3 Gnd 1.32fF
C1687 AND4Bit_0/AND2IN_1/NOT_0/in Gnd 0.37fF
C1688 AND4Bit_0/AND2IN_1/NOT_0/w_n7_n3# Gnd 0.61fF
C1689 AND4Bit_0/AND2IN_1/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1690 OR3IN_0/vin3 Gnd 0.37fF
C1691 AND4Bit_0/AND2IN_0/NOT_0/in Gnd 0.37fF
C1692 AND4Bit_0/AND2IN_0/NOT_0/w_n7_n3# Gnd 0.61fF
C1693 AND4Bit_0/AND2IN_0/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1694 Comparator_0/OR4IN_0/w_n19_n9# Gnd 1.95fF
C1695 Comparator_0/OR4IN_0/vout Gnd 0.71fF
C1696 Comparator_0/OR4IN_0/NOT_0/in Gnd 0.51fF
C1697 Comparator_0/OR4IN_0/NOT_0/w_n7_n3# Gnd 0.61fF
C1698 Comparator_0/NOT_4/w_n7_n3# Gnd 0.61fF
C1699 Comparator_0/NOT_4/out Gnd 22.68fF
C1700 Comparator_0/AND4IN_1/w_n14_n10# Gnd 2.83fF
C1701 Comparator_0/OR4IN_0/vin3 Gnd 1.61fF
C1702 Comparator_0/AND4IN_1/NOT_0/in Gnd 0.45fF
C1703 Comparator_0/AND4IN_1/NOT_0/w_n7_n3# Gnd 0.61fF
C1704 Comparator_0/NOT_3/out Gnd 0.56fF
C1705 Comparator_0/NOT_3/w_n7_n3# Gnd 0.61fF
C1706 Comparator_0/AND4IN_0/w_n14_n10# Gnd 2.83fF
C1707 Comparator_0/AND4IN_0/vout Gnd 0.68fF
C1708 Comparator_0/AND4IN_0/NOT_0/in Gnd 0.45fF
C1709 Comparator_0/AND4IN_0/NOT_0/w_n7_n3# Gnd 0.61fF
C1710 Comparator_0/NOT_2/out Gnd 0.42fF
C1711 Comparator_0/NOT_2/w_n7_n3# Gnd 0.61fF
C1712 Comparator_0/NOT_0/w_n7_n3# Gnd 0.61fF
C1713 Comparator_0/NOT_1/out Gnd 0.43fF
C1714 Comparator_0/NOT_1/w_n7_n3# Gnd 0.61fF
C1715 Comparator_0/AND2IN_3/NOT_0/in Gnd 0.37fF
C1716 Comparator_0/AND2IN_3/NOT_0/w_n7_n3# Gnd 0.61fF
C1717 Comparator_0/NOR2IN_0/vout Gnd 0.03fF
C1718 Comparator_0/AND2IN_3/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1719 Comparator_0/NOT_6/out Gnd 1.41fF
C1720 Comparator_0/AND5IN_0/w_n26_1# Gnd 1.65fF
C1721 Comparator_0/OR4IN_0/vin4 Gnd 1.86fF
C1722 Comparator_0/AND5IN_0/NOT_0/in Gnd 0.65fF
C1723 Comparator_0/AND5IN_0/NOT_0/w_n7_n3# Gnd 0.61fF
C1724 OR3IN_2/vin2 Gnd 2.29fF
C1725 Comparator_0/AND2IN_2/NOT_0/in Gnd 0.37fF
C1726 Comparator_0/AND2IN_2/NOT_0/w_n7_n3# Gnd 0.61fF
C1727 Comparator_0/AND2IN_2/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1728 OR3IN_0/vin2 Gnd 1.28fF
C1729 Comparator_0/AND2IN_1/NOT_0/in Gnd 0.37fF
C1730 Comparator_0/AND2IN_1/NOT_0/w_n7_n3# Gnd 0.61fF
C1731 Comparator_0/AND2IN_1/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1732 Comparator_0/AND2IN_0/NOT_0/in Gnd 0.37fF
C1733 Comparator_0/AND2IN_0/NOT_0/w_n7_n3# Gnd 0.61fF
C1734 Comparator_0/AND2IN_0/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1735 Comparator_0/NOR2IN_0/w_n19_n9# Gnd 1.37fF
C1736 Comparator_0/NOT_5/in Gnd 4.73fF
C1737 Comparator_0/XOR2IN_3/NAND2IN_3/vin1 Gnd 0.54fF
C1738 Comparator_0/XOR2IN_3/NAND2IN_3/w_n16_n4# Gnd 1.16fF
C1739 Comparator_0/XOR2IN_3/NAND2IN_3/vin2 Gnd 0.55fF
C1740 Comparator_0/XOR2IN_3/NAND2IN_2/vin2 Gnd 0.80fF
C1741 Comparator_0/XOR2IN_3/NAND2IN_2/w_n16_n4# Gnd 1.16fF
C1742 Comparator_0/XOR2IN_3/NAND2IN_1/w_n16_n4# Gnd 1.16fF
C1743 Enable_1/voutb3 Gnd 12.65fF
C1744 Enable_1/vouta3 Gnd 2.82fF
C1745 Comparator_0/XOR2IN_3/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1746 Comparator_0/NOT_4/in Gnd 0.67fF
C1747 Comparator_0/XOR2IN_2/NAND2IN_3/vin1 Gnd 0.54fF
C1748 Comparator_0/XOR2IN_2/NAND2IN_3/w_n16_n4# Gnd 1.16fF
C1749 Comparator_0/XOR2IN_2/NAND2IN_3/vin2 Gnd 0.55fF
C1750 Comparator_0/XOR2IN_2/NAND2IN_2/vin2 Gnd 0.80fF
C1751 Comparator_0/XOR2IN_2/NAND2IN_2/w_n16_n4# Gnd 1.16fF
C1752 Comparator_0/XOR2IN_2/NAND2IN_1/w_n16_n4# Gnd 1.16fF
C1753 Enable_1/voutb2 Gnd 2.64fF
C1754 Enable_1/vouta2 Gnd 3.53fF
C1755 Comparator_0/XOR2IN_2/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1756 Comparator_0/NOT_6/in Gnd 0.86fF
C1757 Comparator_0/XOR2IN_1/NAND2IN_3/vin1 Gnd 0.54fF
C1758 Comparator_0/XOR2IN_1/NAND2IN_3/w_n16_n4# Gnd 1.16fF
C1759 Comparator_0/XOR2IN_1/NAND2IN_3/vin2 Gnd 0.55fF
C1760 Comparator_0/XOR2IN_1/NAND2IN_2/vin2 Gnd 0.80fF
C1761 Comparator_0/XOR2IN_1/NAND2IN_2/w_n16_n4# Gnd 1.16fF
C1762 Comparator_0/XOR2IN_1/NAND2IN_1/w_n16_n4# Gnd 1.16fF
C1763 Enable_1/vouta1 Gnd 11.15fF
C1764 Comparator_0/XOR2IN_1/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1765 Comparator_0/XOR2IN_0/NAND2IN_3/vin1 Gnd 0.54fF
C1766 Comparator_0/XOR2IN_0/NAND2IN_3/w_n16_n4# Gnd 1.16fF
C1767 Comparator_0/XOR2IN_0/NAND2IN_3/vin2 Gnd 0.55fF
C1768 Comparator_0/XOR2IN_0/NAND2IN_2/vin2 Gnd 0.80fF
C1769 Comparator_0/XOR2IN_0/NAND2IN_2/w_n16_n4# Gnd 1.16fF
C1770 Comparator_0/XOR2IN_0/NAND2IN_1/w_n16_n4# Gnd 1.16fF
C1771 Enable_1/vouta0 Gnd 3.93fF
C1772 Comparator_0/XOR2IN_0/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1773 Comparator_0/NOT_5/out Gnd 1.69fF
C1774 Comparator_0/AND3IN_0/w_n14_n10# Gnd 2.32fF
C1775 Comparator_0/OR4IN_0/vin2 Gnd 1.19fF
C1776 Comparator_0/AND3IN_0/NOT_0/in Gnd 0.44fF
C1777 Comparator_0/AND3IN_0/NOT_0/w_n7_n3# Gnd 0.61fF
C1778 Comparator_0/NOT_7/out Gnd 0.42fF
C1779 Comparator_0/NOT_7/w_n7_n3# Gnd 0.61fF
C1780 Comparator_0/NOT_6/w_n7_n3# Gnd 0.61fF
C1781 Comparator_0/NOT_5/w_n7_n3# Gnd 0.61fF
C1782 OR2IN_1/w_n19_n9# Gnd 1.40fF
C1783 OR2IN_1/NOT_0/in Gnd 0.42fF
C1784 OR2IN_1/NOT_0/w_n7_n3# Gnd 0.61fF
C1785 OR2IN_0/w_n19_n9# Gnd 1.40fF
C1786 OR2IN_0/NOT_0/in Gnd 0.42fF
C1787 OR2IN_0/NOT_0/w_n7_n3# Gnd 0.61fF
C1788 OR3IN_2/w_n19_n9# Gnd 1.71fF
C1789 OR3IN_2/NOT_0/in Gnd 0.45fF
C1790 OR3IN_2/NOT_0/w_n7_n3# Gnd 0.61fF
C1791 OR3IN_1/w_n19_n9# Gnd 1.71fF
C1792 vout1 Gnd 0.09fF
C1793 OR3IN_1/NOT_0/in Gnd 0.45fF
C1794 OR3IN_1/NOT_0/w_n7_n3# Gnd 0.61fF
C1795 OR3IN_0/w_n19_n9# Gnd 1.71fF
C1796 vout0 Gnd 0.10fF
C1797 OR3IN_0/NOT_0/in Gnd 0.45fF
C1798 OR3IN_0/NOT_0/w_n7_n3# Gnd 0.61fF
C1799 Decoder_0/NOT_0/w_n7_n3# Gnd 0.61fF
C1800 Decoder_0/NOT_1/w_n7_n3# Gnd 0.61fF
C1801 Decoder_0/AND4Bit_0/AND2IN_3/NOT_0/in Gnd 0.37fF
C1802 Decoder_0/AND4Bit_0/AND2IN_3/NOT_0/w_n7_n3# Gnd 0.61fF
C1803 Decoder_0/AND4Bit_0/AND2IN_3/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1804 Decoder_0/AND4Bit_0/AND2IN_2/NOT_0/in Gnd 0.37fF
C1805 Decoder_0/AND4Bit_0/AND2IN_2/NOT_0/w_n7_n3# Gnd 0.61fF
C1806 vinSel1 Gnd 1.24fF
C1807 Decoder_0/AND4Bit_0/AND2IN_2/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1808 Decoder_0/AND4Bit_0/AND2IN_1/NOT_0/in Gnd 0.37fF
C1809 Decoder_0/AND4Bit_0/AND2IN_1/NOT_0/w_n7_n3# Gnd 0.61fF
C1810 vinSel0 Gnd 1.05fF
C1811 Decoder_0/AND4Bit_0/AND2IN_1/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C1812 OR2IN_0/vin1 Gnd 0.46fF
C1813 Decoder_0/AND4Bit_0/AND2IN_0/NOT_0/in Gnd 0.37fF
C1814 Decoder_0/AND4Bit_0/AND2IN_0/NOT_0/w_n7_n3# Gnd 0.61fF
C1815 Decoder_0/NOT_0/out Gnd 0.94fF
C1816 Decoder_0/NOT_1/out Gnd 2.59fF
C1817 Decoder_0/AND4Bit_0/AND2IN_0/NAND2IN_0/w_n16_n4# Gnd 1.16fF

.tran 1n 200n

.measure tran trise 
+ TRIG v(vinb3) VAL = 'SUPPLY/2' RISE =1
+ TARG v(vout2) VAL = 'SUPPLY/2' RISE =1 

.measure tran tfall 
+ TRIG v(vinb3) VAL = 'SUPPLY/2' FALL =1 
+ TARG v(vout2) VAL = 'SUPPLY/2' FALL=1

.measure tran tpd param = '(trise + tfall)/2' goal = 0
        

.control
run
quit
.end
.endc