* SPICE3 file created from fullAdder.ext - technology: scmos

.option scale=0.09u
.include TSMC_180nm.txt

.param SUPPLY = 1.8
.global gnd

Vdd vdd gnd 'SUPPLY'

V_in_3 vcin gnd PULSE(1.8 0 0ns 100ps 100ps 80ns 160ns)
V_in_2 vin2 gnd PULSE(1.8 0 0ns 100ps 100ps 40ns 80ns)
V_in_1 vin1 gnd PULSE(1.8 0 0ns 100ps 100ps 20ns 40ns)


M1000 XOR2IN_0/NAND2IN_0/a_n1_n23# vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=300 ps=270
M1001 XOR2IN_0/NAND2IN_2/vin2 vin1 vdd XOR2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=562 ps=462
M1002 XOR2IN_0/NAND2IN_2/vin2 vin2 XOR2IN_0/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1003 XOR2IN_0/NAND2IN_2/vin2 vin2 vdd XOR2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 XOR2IN_0/NAND2IN_1/a_n1_n23# vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1005 XOR2IN_0/NAND2IN_3/vin1 vin1 vdd XOR2IN_0/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1006 XOR2IN_0/NAND2IN_3/vin1 XOR2IN_0/NAND2IN_2/vin2 XOR2IN_0/NAND2IN_1/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1007 XOR2IN_0/NAND2IN_3/vin1 XOR2IN_0/NAND2IN_2/vin2 vdd XOR2IN_0/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 XOR2IN_0/NAND2IN_2/a_n1_n23# vin2 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1009 XOR2IN_0/NAND2IN_3/vin2 vin2 vdd XOR2IN_0/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1010 XOR2IN_0/NAND2IN_3/vin2 XOR2IN_0/NAND2IN_2/vin2 XOR2IN_0/NAND2IN_2/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1011 XOR2IN_0/NAND2IN_3/vin2 XOR2IN_0/NAND2IN_2/vin2 vdd XOR2IN_0/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1012 XOR2IN_0/NAND2IN_3/a_n1_n23# XOR2IN_0/NAND2IN_3/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1013 XOR2IN_1/vin1 XOR2IN_0/NAND2IN_3/vin1 vdd XOR2IN_0/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1014 XOR2IN_1/vin1 XOR2IN_0/NAND2IN_3/vin2 XOR2IN_0/NAND2IN_3/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1015 XOR2IN_1/vin1 XOR2IN_0/NAND2IN_3/vin2 vdd XOR2IN_0/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1016 XOR2IN_1/NAND2IN_0/a_n1_n23# XOR2IN_1/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1017 XOR2IN_1/NAND2IN_2/vin2 XOR2IN_1/vin1 vdd XOR2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1018 XOR2IN_1/NAND2IN_2/vin2 vcin XOR2IN_1/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1019 XOR2IN_1/NAND2IN_2/vin2 vcin vdd XOR2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1020 XOR2IN_1/NAND2IN_1/a_n1_n23# XOR2IN_1/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1021 XOR2IN_1/NAND2IN_3/vin1 XOR2IN_1/vin1 vdd XOR2IN_1/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1022 XOR2IN_1/NAND2IN_3/vin1 XOR2IN_1/NAND2IN_2/vin2 XOR2IN_1/NAND2IN_1/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1023 XOR2IN_1/NAND2IN_3/vin1 XOR2IN_1/NAND2IN_2/vin2 vdd XOR2IN_1/NAND2IN_1/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1024 XOR2IN_1/NAND2IN_2/a_n1_n23# vcin gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1025 XOR2IN_1/NAND2IN_3/vin2 vcin vdd XOR2IN_1/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1026 XOR2IN_1/NAND2IN_3/vin2 XOR2IN_1/NAND2IN_2/vin2 XOR2IN_1/NAND2IN_2/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1027 XOR2IN_1/NAND2IN_3/vin2 XOR2IN_1/NAND2IN_2/vin2 vdd XOR2IN_1/NAND2IN_2/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1028 XOR2IN_1/NAND2IN_3/a_n1_n23# XOR2IN_1/NAND2IN_3/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1029 vout XOR2IN_1/NAND2IN_3/vin1 vdd XOR2IN_1/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1030 vout XOR2IN_1/NAND2IN_3/vin2 XOR2IN_1/NAND2IN_3/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1031 vout XOR2IN_1/NAND2IN_3/vin2 vdd XOR2IN_1/NAND2IN_3/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1032 AND2IN_0/NAND2IN_0/a_n1_n23# vin1 gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1033 AND2IN_0/NOT_0/in vin1 vdd AND2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1034 AND2IN_0/NOT_0/in vin2 AND2IN_0/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1035 AND2IN_0/NOT_0/in vin2 vdd AND2IN_0/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1036 OR2IN_0/vin2 AND2IN_0/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1037 OR2IN_0/vin2 AND2IN_0/NOT_0/in vdd AND2IN_0/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1038 vcout OR2IN_0/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1039 vcout OR2IN_0/NOT_0/in vdd OR2IN_0/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1040 OR2IN_0/NOT_0/in OR2IN_0/vin2 OR2IN_0/a_0_1# OR2IN_0/w_n19_n9# CMOSP w=12 l=2
+  ad=72 pd=36 as=48 ps=32
M1041 OR2IN_0/NOT_0/in OR2IN_0/vin2 gnd Gnd CMOSN w=4 l=2
+  ad=60 pd=46 as=0 ps=0
M1042 OR2IN_0/a_0_1# OR2IN_0/vin1 vdd OR2IN_0/w_n19_n9# CMOSP w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1043 OR2IN_0/NOT_0/in OR2IN_0/vin1 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1044 AND2IN_1/NAND2IN_0/a_n1_n23# vcin gnd Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1045 AND2IN_1/NOT_0/in vcin vdd AND2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1046 AND2IN_1/NOT_0/in XOR2IN_1/vin1 AND2IN_1/NAND2IN_0/a_n1_n23# Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1047 AND2IN_1/NOT_0/in XOR2IN_1/vin1 vdd AND2IN_1/NAND2IN_0/w_n16_n4# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1048 OR2IN_0/vin1 AND2IN_1/NOT_0/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1049 OR2IN_0/vin1 AND2IN_1/NOT_0/in vdd AND2IN_1/NOT_0/w_n7_n3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
C0 XOR2IN_1/NAND2IN_3/vin1 XOR2IN_1/NAND2IN_2/vin2 0.06fF
C1 vdd OR2IN_0/vin2 0.06fF
C2 vcin gnd 0.40fF
C3 OR2IN_0/w_n19_n9# OR2IN_0/NOT_0/in 0.05fF
C4 vin2 AND2IN_0/NOT_0/in 0.06fF
C5 XOR2IN_1/NAND2IN_3/w_n16_n4# vout 0.08fF
C6 XOR2IN_0/NAND2IN_1/w_n16_n4# vin1 0.10fF
C7 vcin OR2IN_0/vin2 0.06fF
C8 XOR2IN_0/NAND2IN_0/w_n16_n4# XOR2IN_0/NAND2IN_2/vin2 0.08fF
C9 vdd AND2IN_0/NAND2IN_0/w_n16_n4# 0.11fF
C10 AND2IN_1/NAND2IN_0/w_n16_n4# XOR2IN_1/vin1 0.10fF
C11 gnd OR2IN_0/NOT_0/in 0.11fF
C12 XOR2IN_1/vin1 XOR2IN_1/NAND2IN_1/w_n16_n4# 0.10fF
C13 vdd XOR2IN_1/NAND2IN_2/w_n16_n4# 0.11fF
C14 XOR2IN_0/NAND2IN_3/vin1 gnd 0.06fF
C15 OR2IN_0/vin2 OR2IN_0/NOT_0/in 0.08fF
C16 XOR2IN_1/NAND2IN_3/w_n16_n4# XOR2IN_1/NAND2IN_3/vin2 0.10fF
C17 XOR2IN_0/NAND2IN_3/vin2 XOR2IN_0/NAND2IN_2/vin2 0.06fF
C18 vdd XOR2IN_0/NAND2IN_2/w_n16_n4# 0.11fF
C19 XOR2IN_1/NAND2IN_0/w_n16_n4# XOR2IN_1/NAND2IN_2/vin2 0.08fF
C20 vdd vcin 0.06fF
C21 vcin XOR2IN_1/NAND2IN_2/w_n16_n4# 0.10fF
C22 gnd XOR2IN_0/NAND2IN_2/vin2 0.19fF
C23 vdd vout 0.08fF
C24 XOR2IN_0/NAND2IN_1/w_n16_n4# vdd 0.11fF
C25 vin2 XOR2IN_0/NAND2IN_0/w_n16_n4# 0.10fF
C26 gnd XOR2IN_1/NAND2IN_2/vin2 0.19fF
C27 vdd XOR2IN_0/NAND2IN_3/vin1 0.43fF
C28 XOR2IN_1/vin1 AND2IN_1/NOT_0/in 0.06fF
C29 vdd XOR2IN_1/NAND2IN_3/vin2 0.08fF
C30 AND2IN_1/NAND2IN_0/w_n16_n4# vdd 0.14fF
C31 AND2IN_0/NOT_0/w_n7_n3# AND2IN_0/NOT_0/in 0.07fF
C32 XOR2IN_1/NAND2IN_3/vin2 XOR2IN_1/NAND2IN_2/w_n16_n4# 0.08fF
C33 vin1 vin2 0.27fF
C34 vdd XOR2IN_1/NAND2IN_1/w_n16_n4# 0.11fF
C35 vdd XOR2IN_0/NAND2IN_2/vin2 0.15fF
C36 vdd AND2IN_1/NOT_0/w_n7_n3# 0.06fF
C37 vin2 gnd 0.21fF
C38 XOR2IN_0/NAND2IN_2/w_n16_n4# XOR2IN_0/NAND2IN_2/vin2 0.10fF
C39 AND2IN_1/NOT_0/in gnd 0.05fF
C40 AND2IN_1/NAND2IN_0/w_n16_n4# vcin 0.10fF
C41 vdd XOR2IN_1/NAND2IN_2/vin2 0.08fF
C42 XOR2IN_1/NAND2IN_2/w_n16_n4# XOR2IN_1/NAND2IN_2/vin2 0.10fF
C43 XOR2IN_0/NAND2IN_1/w_n16_n4# XOR2IN_0/NAND2IN_3/vin1 0.08fF
C44 vout XOR2IN_1/NAND2IN_3/vin2 0.06fF
C45 OR2IN_0/vin1 OR2IN_0/w_n19_n9# 0.16fF
C46 AND2IN_0/NOT_0/in gnd 0.05fF
C47 XOR2IN_1/vin1 XOR2IN_0/NAND2IN_3/w_n16_n4# 0.08fF
C48 vcin XOR2IN_1/NAND2IN_2/vin2 0.39fF
C49 XOR2IN_0/NAND2IN_3/vin2 XOR2IN_0/NAND2IN_3/w_n16_n4# 0.10fF
C50 XOR2IN_0/NAND2IN_1/w_n16_n4# XOR2IN_0/NAND2IN_2/vin2 0.10fF
C51 vin2 AND2IN_0/NAND2IN_0/w_n16_n4# 0.10fF
C52 OR2IN_0/vin1 gnd 0.26fF
C53 OR2IN_0/NOT_0/w_n7_n3# vcout 0.03fF
C54 XOR2IN_1/NAND2IN_3/w_n16_n4# XOR2IN_1/NAND2IN_3/vin1 0.10fF
C55 vdd vin2 0.12fF
C56 XOR2IN_0/NAND2IN_3/vin1 XOR2IN_0/NAND2IN_2/vin2 0.06fF
C57 XOR2IN_1/NAND2IN_3/vin1 gnd 0.06fF
C58 vdd AND2IN_1/NOT_0/in 0.08fF
C59 OR2IN_0/vin1 OR2IN_0/vin2 0.11fF
C60 vin2 XOR2IN_0/NAND2IN_2/w_n16_n4# 0.10fF
C61 AND2IN_0/NAND2IN_0/w_n16_n4# AND2IN_0/NOT_0/in 0.08fF
C62 vdd AND2IN_0/NOT_0/in 0.08fF
C63 XOR2IN_1/vin1 XOR2IN_1/NAND2IN_0/w_n16_n4# 0.10fF
C64 XOR2IN_1/NAND2IN_3/vin2 XOR2IN_1/NAND2IN_2/vin2 0.06fF
C65 vin1 XOR2IN_0/NAND2IN_0/w_n16_n4# 0.10fF
C66 XOR2IN_1/vin1 XOR2IN_0/NAND2IN_3/vin2 0.06fF
C67 XOR2IN_1/NAND2IN_1/w_n16_n4# XOR2IN_1/NAND2IN_2/vin2 0.10fF
C68 OR2IN_0/vin1 vdd 0.06fF
C69 OR2IN_0/NOT_0/w_n7_n3# vdd 0.06fF
C70 vdd XOR2IN_1/NAND2IN_3/vin1 0.43fF
C71 XOR2IN_1/vin1 gnd 0.52fF
C72 vdd XOR2IN_0/NAND2IN_3/w_n16_n4# 0.11fF
C73 AND2IN_0/NOT_0/w_n7_n3# OR2IN_0/vin2 0.03fF
C74 vin1 gnd 0.40fF
C75 AND2IN_1/NAND2IN_0/w_n16_n4# AND2IN_1/NOT_0/in 0.08fF
C76 vcout gnd 0.07fF
C77 vin2 XOR2IN_0/NAND2IN_2/vin2 0.39fF
C78 OR2IN_0/w_n19_n9# OR2IN_0/vin2 0.12fF
C79 AND2IN_1/NOT_0/in AND2IN_1/NOT_0/w_n7_n3# 0.07fF
C80 OR2IN_0/NOT_0/w_n7_n3# OR2IN_0/NOT_0/in 0.07fF
C81 vdd XOR2IN_0/NAND2IN_0/w_n16_n4# 0.11fF
C82 vdd AND2IN_0/NOT_0/w_n7_n3# 0.09fF
C83 OR2IN_0/vin2 gnd 0.27fF
C84 vdd XOR2IN_1/NAND2IN_0/w_n16_n4# 0.11fF
C85 XOR2IN_1/vin1 vdd 0.21fF
C86 XOR2IN_0/NAND2IN_3/w_n16_n4# XOR2IN_0/NAND2IN_3/vin1 0.10fF
C87 vdd XOR2IN_0/NAND2IN_3/vin2 0.08fF
C88 vin1 AND2IN_0/NAND2IN_0/w_n16_n4# 0.10fF
C89 vdd OR2IN_0/w_n19_n9# 0.09fF
C90 XOR2IN_0/NAND2IN_3/vin2 XOR2IN_0/NAND2IN_2/w_n16_n4# 0.08fF
C91 OR2IN_0/vin1 AND2IN_1/NOT_0/w_n7_n3# 0.03fF
C92 vcin XOR2IN_1/NAND2IN_0/w_n16_n4# 0.10fF
C93 vdd vin1 0.06fF
C94 XOR2IN_1/vin1 vcin 0.26fF
C95 XOR2IN_1/NAND2IN_3/w_n16_n4# vdd 0.11fF
C96 vdd vcout 0.06fF
C97 XOR2IN_1/NAND2IN_1/w_n16_n4# XOR2IN_1/NAND2IN_3/vin1 0.08fF
C98 vdd gnd 0.39fF
C99 gnd Gnd 0.01fF
C100 AND2IN_1/NOT_0/in Gnd 0.37fF
C101 AND2IN_1/NOT_0/w_n7_n3# Gnd 0.61fF
C102 AND2IN_1/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C103 OR2IN_0/w_n19_n9# Gnd 1.40fF
C104 vcout Gnd 0.09fF
C105 OR2IN_0/NOT_0/in Gnd 0.42fF
C106 OR2IN_0/NOT_0/w_n7_n3# Gnd 0.61fF
C107 vdd Gnd 3.50fF
C108 AND2IN_0/NOT_0/in Gnd 0.37fF
C109 AND2IN_0/NOT_0/w_n7_n3# Gnd 0.61fF
C110 AND2IN_0/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C111 vout Gnd 0.22fF
C112 XOR2IN_1/NAND2IN_3/vin1 Gnd 0.54fF
C113 XOR2IN_1/NAND2IN_3/w_n16_n4# Gnd 1.16fF
C114 XOR2IN_1/NAND2IN_3/vin2 Gnd 0.55fF
C115 XOR2IN_1/NAND2IN_2/vin2 Gnd 0.80fF
C116 XOR2IN_1/NAND2IN_2/w_n16_n4# Gnd 1.16fF
C117 XOR2IN_1/NAND2IN_1/w_n16_n4# Gnd 1.16fF
C118 vcin Gnd 6.53fF
C119 XOR2IN_1/vin1 Gnd 3.73fF
C120 XOR2IN_1/NAND2IN_0/w_n16_n4# Gnd 1.16fF
C121 XOR2IN_0/NAND2IN_3/vin1 Gnd 0.54fF
C122 XOR2IN_0/NAND2IN_3/w_n16_n4# Gnd 1.16fF
C123 XOR2IN_0/NAND2IN_3/vin2 Gnd 0.55fF
C124 XOR2IN_0/NAND2IN_2/vin2 Gnd 0.80fF
C125 XOR2IN_0/NAND2IN_2/w_n16_n4# Gnd 1.16fF
C126 XOR2IN_0/NAND2IN_1/w_n16_n4# Gnd 1.16fF
C127 vin2 Gnd 2.21fF
C128 vin1 Gnd 5.54fF
C129 XOR2IN_0/NAND2IN_0/w_n16_n4# Gnd 1.16fF

.tran 1n 160n

.control
run

set color0 = rgb:f/f/e
set color1 = black
plot v(vin1) v(vin2)+2 v(vcin)+4 v(vout)+6 v(vcout)+8

hardcopy image.ps v(vin1) v(vin2)+2 v(vcin)+4 v(vout)+6 v(vcout)+8
.end
.endc