* SPICE3 file created from NOR2IN.ext - technology: scmos

.include TSMC_180nm.txt
.option scale=0.09u

.param SUPPLY = 1.8
.global gnd

Vdd vdd gnd 'SUPPLY'

V_in_a vin1 gnd PULSE(1.8 0 0ns 100ps 100ps 20ns 40ns)
V_in_b vin2 gnd PULSE(1.8 0 0ns 100ps 100ps 40ns 80ns)

M1000 vout vin2 a_0_1# w_n19_n9# CMOSP w=12 l=2
+  ad=72 pd=36 as=48 ps=32
M1001 vout vin2 gnd Gnd CMOSN w=4 l=2
+  ad=60 pd=46 as=40 ps=36
M1002 a_0_1# vin1 vdd w_n19_n9# CMOSP w=12 l=2
+  ad=0 pd=0 as=72 ps=36
M1003 vout vin1 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
C0 w_n19_n9# vdd 0.09fF
C1 vin2 vin1 0.11fF
C2 vout gnd 0.11fF
C3 w_n19_n9# vout 0.05fF
C4 vin2 vout 0.08fF
C5 vin1 gnd 0.12fF
C6 w_n19_n9# vin2 0.12fF
C7 w_n19_n9# vin1 0.16fF
C8 gnd Gnd 0.15fF
C9 vout Gnd 0.17fF
C10 vdd Gnd 0.07fF
C11 vin2 Gnd 0.26fF
C12 vin1 Gnd 0.32fF
C13 w_n19_n9# Gnd 1.37fF

.tran 1n 80n

.control
run
set color0 = rgb:f/f/e
set color1 = black
plot v(vin1) v(vin2)+2 (vout)+4
hardcopy image.ps v(vin1) v(vin2)+2 (vout)+4
.end
.endc