magic
tech scmos
timestamp 1698770891
<< metal1 >>
rect 74 206 80 209
rect 233 206 310 209
rect 307 131 310 206
rect 301 106 312 109
rect 331 105 342 108
rect 308 89 317 92
rect 80 71 83 85
rect -23 57 -14 60
rect -23 0 -14 3
<< m2contact >>
rect 303 87 308 92
<< metal2 >>
rect 219 7 222 100
rect 303 7 306 87
rect 219 4 306 7
use NOT  NOT_0
timestamp 1698475750
transform 1 0 314 0 1 115
box -7 -26 25 19
use XOR2IN  XOR2IN_0
timestamp 1698769192
transform 1 0 91 0 1 108
box -106 -118 213 101
<< labels >>
rlabel metal1 75 207 76 208 5 vdd
rlabel metal1 81 75 82 76 1 gnd
rlabel metal1 -21 58 -20 59 3 vin1
rlabel metal1 -22 1 -21 2 3 vin2
rlabel metal1 339 106 340 107 7 vout
<< end >>
