Absolute value using 4bitAdder

.include TSMC_180nm.txt
.include All_Gates.sub

.subckt fullAdder Cout S A B Cin vdd gnd
    X1 S1out A B vdd gnd XOR2IN
    X2 S S1out Cin vdd gnd XOR2IN
    X3 C1out A B vdd gnd AND2IN
    X4 C2out S1out Cin vdd gnd AND2IN
    X5 Cout C1out C2out vdd gnd OR2IN
.ends fullAdder

.subckt 4bitAdder s3 s2 s1 s0 Carry node_a3 node_a2 node_a1 node_a0 node_b3 node_b2 node_b1 node_b0 node_m vdd gnd
    X1 B0 node_m node_b0 vdd gnd XOR2IN
    X2 B1 node_m node_b1 vdd gnd XOR2IN
    X3 B2 node_m node_b2 vdd gnd XOR2IN
    X4 B3 node_m node_b3 vdd gnd XOR2IN
    X5 Cout0 s0 node_a0 B0 node_m vdd gnd fullAdder
    X6 Cout1 s1 node_a1 B1 Cout0 vdd gnd fullAdder
    X7 Cout2 s2 node_a2 B2 Cout1 vdd gnd fullAdder
    X8 Carry s3 node_a3 B3 Cout2 vdd gnd fullAdder
.ends 4bitAdder 

.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd vdd gnd 'SUPPLY'

V_in_a3 node_a3 gnd DC 0
V_in_a2 node_a2 gnd DC 0
V_in_a1 node_a1 gnd DC 0
V_in_a0 node_a0 gnd DC 0

V_in_b3 node_b3 gnd PULSE(0 1.8 0ns 100ps 100ps 160ns 320ns)
V_in_b2 node_b2 gnd PULSE(0 1.8 0ns 100ps 100ps 80ns 160ns)
V_in_b1 node_b1 gnd PULSE(0 1.8 0ns 100ps 100ps 40ns 80ns)
V_in_b0 node_b0 gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)


X_add node_out3 node_out2 node_out1 node_out0 Carry node_a3 node_a2 node_a1 node_a0 node_b3 node_b2 node_b1 node_b0 node_b3 vdd gnd 4bitAdder

C1 node_out0 gnd 100f
C2 node_out1 gnd 100f
C3 node_out2 gnd 100f
C4 node_out3 gnd 100f

.tran 1n 320n

.control
run

set color0 = rgb:f/f/e
set color1 = black
plot v(node_b0) v(node_out0)+8 v(node_b1)+2 v(node_out1)+10 v(node_b2)+4 v(node_out2)+12 v(node_b3)+6 v(node_out3)+14

hardcopy image.ps v(node_b0) v(node_out0)+8 v(node_b1)+2 v(node_out1)+10 v(node_b2)+4 v(node_out2)+12 v(node_b3)+6 v(node_out3)+14
.end
.endc



