Question No 2 Ring Oscillator

.include TSMC_180nm.txt
.include All_Gates.sub

.subckt RingOscillator Out vdd gnd
    X1 o1 Out vdd gnd NOT
    X2 o2 o1 vdd gnd NOT
    X3 Out o2 vdd gnd NOT
.ends RingOscillator

.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd vdd gnd 'SUPPLY'

.ic V(Out)= 0V
Xr Out vdd gnd RingOscillator
* Xn Out Out vdd gnd NOT

C1 Out gnd 50f

.tran 1n 20n

.control
run

set color0 = rgb:f/f/e
set color1 = black
plot v(Out)
hardcopy image.ps v(Out)
.end
.endc
