magic
tech scmos
timestamp 1698684844
<< nwell >>
rect -14 -10 54 24
<< ntransistor >>
rect 0 -30 2 -26
rect 17 -30 19 -26
rect 34 -30 36 -26
<< ptransistor >>
rect 0 8 2 12
rect 17 8 19 12
rect 34 8 36 12
<< ndiffusion >>
rect -1 -30 0 -26
rect 2 -30 17 -26
rect 19 -30 34 -26
rect 36 -30 37 -26
<< pdiffusion >>
rect -1 8 0 12
rect 2 8 3 12
rect 16 8 17 12
rect 19 8 20 12
rect 33 8 34 12
rect 36 8 37 12
<< ndcontact >>
rect -5 -30 -1 -26
rect 37 -30 41 -26
<< pdcontact >>
rect -5 8 -1 12
rect 3 8 7 12
rect 12 8 16 12
rect 20 8 24 12
rect 29 8 33 12
rect 37 8 41 12
<< polysilicon >>
rect 0 12 2 17
rect 17 12 19 17
rect 34 12 36 17
rect 0 -26 2 8
rect 17 -26 19 8
rect 34 -26 36 8
rect 0 -49 2 -30
rect 17 -49 19 -30
rect 34 -49 36 -30
<< polycontact >>
rect -1 -53 3 -49
rect 16 -53 20 -49
rect 33 -53 37 -49
<< metal1 >>
rect -14 24 68 27
rect -5 12 -2 24
rect 12 12 15 24
rect 29 12 32 24
rect 4 -16 7 8
rect 21 -16 24 8
rect 38 -16 41 8
rect 65 6 68 24
rect 4 -19 70 -16
rect 38 -26 41 -19
rect 91 -20 100 -17
rect -18 -30 -5 -26
rect -18 -33 -15 -30
rect -18 -36 85 -33
rect -1 -59 3 -53
rect 16 -59 20 -53
rect 33 -59 37 -53
use NOT  NOT_0
timestamp 1698475750
transform 1 0 72 0 1 -10
box -7 -26 25 19
<< labels >>
rlabel metal1 26 25 27 26 5 vdd
rlabel metal1 -11 -29 -10 -28 1 gnd
rlabel metal1 95 -19 96 -18 7 vout
rlabel metal1 0 -56 1 -55 1 vin1
rlabel metal1 17 -56 18 -55 1 vin2
rlabel metal1 34 -56 35 -55 1 vin3
<< end >>
