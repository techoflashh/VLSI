Question No 3 MajorityFunction

.include TSMC_180nm.txt
.include All_Gates.sub

.subckt MUX Out A3 A2 A1 A0 S1 S0 vdd gnd
    X1 S1c S1 vdd gnd NOT
    X2 S0c S0 vdd gnd NOT
    X3 Out0 A0 S1c S0c vdd gnd AND3IN
    X4 Out1 A1 S1c S0 vdd gnd AND3IN
    X5 Out2 A2 S1 S0c vdd gnd AND3IN
    X6 Out3 A3 S1 S0 vdd gnd AND3IN
    X7 Out Out0 Out1 Out2 Out3 vdd gnd OR4IN
.ends MUX

.subckt MajorityFunction Out A2 A1 A0 vdd gnd
    X1 Out vdd A0 A0 gnd A2 A1 vdd gnd MUX
.ends MajorityFunction

.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd vdd gnd 'SUPPLY'

V_in_a2 node_a2 gnd PULSE(1.8 0 0ns 100ps 100ps 160ns 320ns)
V_in_a1 node_a1 gnd PULSE(1.8 0 0ns 100ps 100ps 80ns 160ns)
V_in_a0 node_a0 gnd PULSE(1.8 0 0ns 100ps 100ps 40ns 80ns)

Xm node_out node_a2 node_a1 node_a0 vdd gnd MajorityFunction 

C1 node_out gnd 50f

.tran 1n 640n

.control
run

set color0 = rgb:f/f/e
set color1 = black
plot v(node_a0) v(node_a1)+2 v(node_a2)+4 v(node_out)+6 
hardcopy image.ps v(node_a0) v(node_a1)+2 v(node_a2)+4 v(node_out)+6 
.end
.endc