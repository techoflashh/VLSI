magic
tech scmos
timestamp 1699694653
<< metal1 >>
rect 705 405 708 427
rect 1496 405 1499 427
rect 2292 405 2295 427
rect -67 389 59 392
rect 617 389 838 392
rect 1357 389 2093 392
rect 2180 389 2440 392
rect -67 -282 -64 389
rect 705 289 708 377
rect 1496 289 1499 374
rect 2292 289 2295 374
rect 3092 289 3095 427
rect -24 240 7 243
rect 736 240 796 243
rect 1532 240 1592 243
rect 2332 240 2392 243
rect -24 -265 -21 240
rect -12 183 6 186
rect -12 -182 -9 183
rect 736 112 739 240
rect 760 183 796 186
rect 760 112 763 183
rect 1532 112 1535 240
rect 1556 183 1592 186
rect 1556 112 1559 183
rect 2332 112 2335 240
rect 2356 183 2392 186
rect 2356 112 2359 183
rect 3146 98 3149 427
rect 694 95 794 98
rect 1496 95 1590 98
rect 2289 95 2390 98
rect 3092 95 3149 98
rect 0 -32 3 25
rect 791 22 794 95
rect 1587 22 1590 95
rect 2387 22 2390 95
rect 32 0 110 3
rect 178 0 891 3
rect 896 0 909 3
rect 965 0 1701 3
rect 1759 0 2495 3
rect 2527 0 3004 3
rect 0 -35 2742 -32
rect 340 -79 343 -35
rect 1107 -103 1110 -35
rect 1933 -115 1936 -35
rect 2739 -101 2742 -35
rect 2739 -104 2769 -101
rect -12 -185 27 -182
rect 340 -269 343 -133
rect 765 -209 795 -206
rect -67 -285 93 -282
rect 244 -285 862 -282
rect 1107 -294 1110 -157
rect 1561 -221 1619 -218
rect -24 -370 -21 -299
rect 1933 -295 1936 -169
rect 2361 -210 2425 -207
rect 736 -305 739 -301
rect -7 -308 739 -305
rect -7 -370 -4 -308
rect 1012 -309 1688 -306
rect 1840 -310 2516 -307
rect 13 -326 1531 -323
rect 13 -370 16 -326
rect 2332 -338 2335 -326
rect 31 -341 2335 -338
rect 31 -370 34 -341
rect 420 -370 423 -353
rect 452 -370 455 -354
rect 478 -370 481 -361
rect 2739 -364 2742 -158
rect 500 -367 2742 -364
rect 2766 -367 2769 -104
rect 500 -370 503 -367
<< m2contact >>
rect 704 400 709 405
rect 1495 400 1500 405
rect 2291 400 2296 405
rect 704 377 709 382
rect 1495 374 1500 379
rect 2291 374 2296 379
rect 735 107 740 112
rect 759 107 764 112
rect 1531 107 1536 112
rect 1555 107 1560 112
rect 2331 107 2336 112
rect 2355 107 2360 112
rect 121 -1 126 4
rect 891 -1 896 4
rect 1715 -1 1720 4
rect 2519 -1 2524 4
rect -25 -270 -20 -265
rect 760 -209 765 -204
rect 339 -274 344 -269
rect 1556 -221 1561 -216
rect -25 -299 -20 -294
rect 735 -301 740 -296
rect 1106 -299 1111 -294
rect 2356 -210 2361 -205
rect 1932 -300 1937 -295
rect 1531 -327 1536 -322
rect 2331 -326 2336 -321
rect 418 -353 423 -348
rect 452 -354 457 -349
rect 478 -361 483 -356
<< metal2 >>
rect 705 382 708 400
rect 1496 379 1499 400
rect 2292 379 2295 400
rect 122 -175 125 -1
rect -24 -294 -21 -270
rect 340 -348 343 -274
rect 736 -296 739 107
rect 760 -204 763 107
rect 892 -199 895 -1
rect 340 -351 418 -348
rect 1107 -349 1110 -299
rect 1532 -322 1535 107
rect 1556 -216 1559 107
rect 1716 -211 1719 -1
rect 457 -352 1110 -349
rect 1933 -356 1936 -300
rect 2332 -321 2335 107
rect 2356 -205 2359 107
rect 2520 -200 2523 -1
rect 483 -359 1936 -356
use fullAdder  fullAdder_0
timestamp 1699609590
transform 1 0 886 0 1 496
box -886 -496 -178 -104
use fullAdder  fullAdder_1
timestamp 1699609590
transform 1 0 1677 0 1 496
box -886 -496 -178 -104
use fullAdder  fullAdder_2
timestamp 1699609590
transform 1 0 2473 0 1 496
box -886 -496 -178 -104
use fullAdder  fullAdder_3
timestamp 1699609590
transform 1 0 3273 0 1 496
box -886 -496 -178 -104
use XOR2IN  XOR2IN_0
timestamp 1698769192
transform -1 0 237 0 -1 -184
box -106 -118 213 101
use XOR2IN  XOR2IN_1
timestamp 1698769192
transform -1 0 1004 0 -1 -208
box -106 -118 213 101
use XOR2IN  XOR2IN_2
timestamp 1698769192
transform -1 0 1830 0 -1 -220
box -106 -118 213 101
use XOR2IN  XOR2IN_3
timestamp 1698769192
transform -1 0 2636 0 -1 -209
box -106 -118 213 101
<< labels >>
rlabel metal1 47 1 48 2 1 gnd
rlabel metal1 -66 -5 -65 -4 3 vdd
rlabel metal1 706 415 707 416 1 vout0
rlabel metal1 1497 412 1498 413 1 vout1
rlabel metal1 2293 412 2294 413 1 vout2
rlabel metal1 3093 405 3094 406 1 vout3
rlabel metal1 3147 405 3148 406 7 vcout
rlabel metal1 -23 -369 -22 -368 1 vina0
rlabel metal1 -6 -369 -5 -368 1 vina1
rlabel metal1 32 -369 33 -368 1 vina3
rlabel metal1 14 -369 15 -368 1 vina2
rlabel metal1 421 -369 422 -368 1 vinb0
rlabel metal1 453 -369 454 -368 1 vinb1
rlabel metal1 479 -369 480 -368 1 vinb2
rlabel metal1 501 -369 502 -368 1 vinb3
rlabel metal1 2767 -366 2768 -365 1 vinM
<< end >>
