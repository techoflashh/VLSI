* SPICE3 file created from not.ext - technology: scmos

.include TSMC_180nm.txt
.option scale=0.09u

.param SUPPLY = 1.8
.global gnd

Vdd vdd gnd 'SUPPLY'

V_in_a in gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)


M1000 out in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=20 ps=18
M1001 out in vdd vdd CMOSP w=5 l=2
+  ad=30 pd=22 as=30 ps=22
C0 vdd vdd 0.06fF
C1 gnd out 0.07fF
C2 in gnd 0.01fF
C3 vdd out 0.03fF
C4 in vdd 0.07fF
C5 out vdd 0.06fF
C6 gnd Gnd 0.06fF
C7 out Gnd 0.05fF
C8 vdd Gnd 0.04fF
C9 in Gnd 0.18fF
C10 vdd Gnd 0.61fF

.tran 1n 800n

.control
run
set color0 = rgb:f/f/e
set color1 = black
plot v(in) v(out)+2
hardcopy image.ps v(in) v(out)+2
.end
.endc
