magic
tech scmos
timestamp 1698495245
<< nwell >>
rect -7 -3 25 16
rect 32 -3 64 16
<< ntransistor >>
rect 8 -19 10 -15
rect -1 -34 1 -30
<< ptransistor >>
rect 8 4 10 9
rect 46 4 48 9
<< ndiffusion >>
rect 7 -19 8 -15
rect 10 -19 12 -15
rect -2 -34 -1 -30
rect 1 -34 3 -30
<< pdiffusion >>
rect 6 4 8 9
rect 10 4 12 9
rect 45 4 46 9
rect 48 4 51 9
<< ndcontact >>
rect 3 -19 7 -15
rect 12 -19 16 -15
rect -6 -34 -2 -30
rect 3 -34 7 -30
<< pdcontact >>
rect 2 4 6 9
rect 12 4 16 9
rect 41 4 45 9
rect 51 4 55 9
<< polysilicon >>
rect 8 9 10 12
rect 46 9 48 12
rect 8 -6 10 4
rect 4 -9 10 -6
rect 8 -15 10 -9
rect 46 -15 48 4
rect 41 -18 48 -15
rect 8 -22 10 -19
rect 46 -27 48 -18
rect -1 -29 48 -27
rect -1 -30 1 -29
rect -1 -37 1 -34
<< polycontact >>
rect 0 -9 4 -5
rect 37 -19 41 -15
<< metal1 >>
rect -7 16 64 19
rect 2 9 5 16
rect 41 9 44 16
rect -3 -9 0 -6
rect 13 -7 16 4
rect 52 -7 55 4
rect 13 -10 55 -7
rect 13 -15 16 -10
rect 32 -18 37 -15
rect 3 -30 6 -19
rect -6 -38 -3 -34
rect -8 -41 -1 -38
<< labels >>
rlabel metal1 6 17 9 18 5 vdd
rlabel metal1 -2 -8 -1 -7 1 vin1
rlabel metal1 33 -17 34 -16 1 vin2
rlabel metal1 25 -9 26 -8 1 vout
rlabel metal1 -5 -40 -4 -39 1 gnd
<< end >>
