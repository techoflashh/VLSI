Question No 5

*temperature

.include TSMC_180nm.txt
.include NAND.sub

.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd vdd gnd 'SUPPLY'

V_in_a nodeA gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)
V_in_b nodeB gnd PULSE(0 1.8 0ns 100ps 100ps 60ns 120ns)

X1 node_out nodeA nodeB vdd gnd NAND

*capacitance

.tran 1n 600n

.measure tran trise
+ TRIG v(nodeA) VAL = 'SUPPLY/2' RISE = 1
+ TARG v(node_out) VAL = 'SUPPLY/2' FALL =1

.measure tran tfall
+ TRIG v(nodeA) VAL = 'SUPPLY/2' FALL = 1
+ TARG v(node_out) VAL = 'SUPPLY/2' RISE =1

.measure tran tpd param = '(trise + tfall)/2' goal = 0 

.control
run

quit
.end
.endc