Testbench for ALU

.include TSMC_180nm.txt
.include ALU.sub

.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd vdd gnd 'SUPPLY'

V_in_a3 node_a3 gnd DC 0
V_in_a2 node_a2 gnd DC 0
V_in_a1 node_a1 gnd DC 0
V_in_a0 node_a0 gnd DC 0

V_in_b3 node_b3 gnd PULSE(0 1.8 0ns 100ps 100ps 60ns 120ns)
V_in_b2 node_b2 gnd PULSE(0 1.8 0ns 100ps 100ps 60ns 120ns)
V_in_b1 node_b1 gnd PULSE(0 1.8 0ns 100ps 100ps 60ns 120ns)
V_in_b0 node_b0 gnd PULSE(0 1.8 0ns 100ps 100ps 60ns 120ns)

V_in_s1 Sel1 gnd DC 0
V_in_s0 Sel0 gnd DC 0

X_ALU CarryOut node_out3 node_out2 node_out1 node_out0 node_a3 node_a2 node_a1 node_a0 node_b3 node_b2 node_b1 node_b0 Sel1 Sel0 vdd gnd ALU


C1 node_out0 gnd 100f
C2 node_out1 gnd 100f
C3 node_out2 gnd 100f
C4 node_out3 gnd 100f
C5 CarryOut gnd 100f

.tran 1n 400n

*targetText

.control
run
quit
.end
.endc