magic
tech scmos
timestamp 1698684672
<< nwell >>
rect -14 -10 69 24
<< ntransistor >>
rect 0 -30 2 -26
rect 17 -30 19 -26
rect 34 -30 36 -26
rect 51 -30 53 -26
<< ptransistor >>
rect 0 8 2 12
rect 17 8 19 12
rect 34 8 36 12
rect 51 8 53 12
<< ndiffusion >>
rect -1 -30 0 -26
rect 2 -30 17 -26
rect 19 -30 34 -26
rect 36 -30 51 -26
rect 53 -30 54 -26
<< pdiffusion >>
rect -1 8 0 12
rect 2 8 3 12
rect 16 8 17 12
rect 19 8 20 12
rect 33 8 34 12
rect 36 8 37 12
rect 50 8 51 12
rect 53 8 54 12
<< ndcontact >>
rect -5 -30 -1 -26
rect 54 -30 58 -26
<< pdcontact >>
rect -5 8 -1 12
rect 3 8 7 12
rect 12 8 16 12
rect 20 8 24 12
rect 29 8 33 12
rect 37 8 41 12
rect 46 8 50 12
rect 54 8 58 12
<< polysilicon >>
rect 0 12 2 17
rect 17 12 19 17
rect 34 12 36 17
rect 51 12 53 17
rect 0 -26 2 8
rect 17 -26 19 8
rect 34 -26 36 8
rect 51 -26 53 8
rect 0 -48 2 -30
rect 17 -48 19 -30
rect 34 -48 36 -30
rect 51 -48 53 -30
<< polycontact >>
rect -1 -52 3 -48
rect 16 -52 20 -48
rect 33 -52 37 -48
rect 50 -52 54 -48
<< metal1 >>
rect -14 24 82 27
rect -5 12 -2 24
rect 12 12 15 24
rect 29 12 32 24
rect 46 12 49 24
rect 4 -16 7 8
rect 21 -16 24 8
rect 38 -16 41 8
rect 55 -16 58 8
rect 79 6 82 24
rect 4 -19 84 -16
rect 55 -26 58 -19
rect 105 -20 114 -17
rect -18 -30 -5 -26
rect -18 -36 -15 -30
rect 75 -36 89 -33
rect -18 -39 78 -36
rect -1 -58 3 -52
rect 16 -58 20 -52
rect 33 -58 37 -52
rect 50 -58 54 -52
use NOT  NOT_0
timestamp 1698475750
transform 1 0 86 0 1 -10
box -7 -26 25 19
<< labels >>
rlabel metal1 26 25 27 26 5 vdd
rlabel metal1 -11 -29 -10 -28 1 gnd
rlabel metal1 109 -19 110 -18 7 vout
rlabel metal1 0 -55 1 -54 1 vin1
rlabel metal1 17 -55 18 -54 1 vin2
rlabel metal1 34 -55 35 -54 1 vin3
rlabel metal1 51 -55 52 -54 1 vin4
<< end >>
