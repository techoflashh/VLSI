magic
tech scmos
timestamp 1699693233
<< metal1 >>
rect 1068 472 1071 515
rect 1137 491 1157 494
rect 1191 491 1308 494
rect 1137 461 1141 491
rect 891 458 913 461
rect 970 458 1141 461
rect 1418 460 1421 522
rect 773 364 815 367
rect 891 364 894 458
rect 1397 457 1421 460
rect 1625 469 1628 522
rect 1625 466 1786 469
rect 1189 447 1268 450
rect 1036 437 1152 440
rect 1001 424 1067 427
rect 1072 424 1120 427
rect 925 387 928 389
rect 944 366 947 392
rect 773 356 776 364
rect 963 359 966 411
rect 985 408 1027 411
rect 1117 406 1120 424
rect 1153 406 1157 414
rect 1117 403 1157 406
rect 1177 402 1181 414
rect 1265 412 1268 447
rect 1383 428 1386 444
rect 1318 412 1321 423
rect 1265 409 1321 412
rect 1625 402 1628 466
rect 1177 399 1628 402
rect 1653 453 1694 456
rect 271 353 658 356
rect 661 353 776 356
rect 271 219 274 353
rect 1030 352 1038 355
rect 1065 352 1180 355
rect 1030 349 1033 352
rect 931 346 1033 349
rect 1653 345 1656 453
rect 1783 419 1786 466
rect 1766 403 1887 406
rect 1722 369 1725 385
rect 1722 366 1874 369
rect 1528 342 1758 345
rect 636 328 660 331
rect 636 282 639 328
rect 679 327 703 330
rect 743 328 749 331
rect 768 327 774 330
rect 944 323 947 328
rect 1028 327 1042 330
rect 1061 326 1069 329
rect 1147 327 1163 330
rect 1182 326 1193 329
rect 937 320 947 323
rect 666 311 811 314
rect 1039 310 1047 313
rect 1055 310 1170 313
rect 922 304 928 307
rect 933 304 962 307
rect 1039 307 1042 310
rect 967 304 1042 307
rect 316 279 639 282
rect 710 279 828 282
rect 316 229 319 279
rect 673 260 736 263
rect 841 263 845 285
rect 1190 284 1193 326
rect 781 260 845 263
rect 858 263 862 284
rect 875 279 1188 282
rect 858 260 1069 263
rect 673 229 676 260
rect 776 241 780 260
rect 1385 250 1405 253
rect 776 238 1459 241
rect 1528 219 1532 342
rect 1871 297 1874 366
rect 1884 284 1887 403
rect 1854 281 2141 284
rect -49 216 95 219
rect 246 216 457 219
rect 603 216 814 219
rect 966 216 1177 219
rect 1328 216 1532 219
rect -49 -81 -46 216
rect 316 116 319 203
rect 673 116 676 203
rect 1033 116 1036 203
rect 1396 116 1399 203
rect 1528 148 1531 216
rect 1753 191 1756 265
rect 1637 188 1756 191
rect 1770 191 1773 266
rect 1788 199 1791 265
rect 1805 209 1808 266
rect 1805 206 2129 209
rect 1788 196 1955 199
rect 1770 188 1793 191
rect 1637 174 1640 188
rect 1615 161 1667 164
rect 1615 140 1618 161
rect 1790 154 1793 188
rect 1808 160 1823 163
rect 1637 117 1640 149
rect 1808 146 1811 160
rect 1952 156 1955 196
rect 1965 170 1983 173
rect 1772 143 1811 146
rect 1965 145 1968 170
rect 1940 142 1968 145
rect 1790 120 1793 131
rect 1772 117 1793 120
rect 1952 119 1955 131
rect 1619 114 1640 117
rect 1934 116 1955 119
rect 2126 118 2129 206
rect 2138 105 2141 281
rect 1660 101 1663 103
rect 1764 101 1816 104
rect 1511 98 1528 101
rect 1607 98 1663 101
rect 1931 100 1981 103
rect 2104 102 2141 105
rect -25 67 3 70
rect 327 67 360 70
rect 687 67 719 70
rect 1050 67 1082 70
rect -25 -64 -22 67
rect 0 -49 3 13
rect 327 -55 330 67
rect 357 -37 360 13
rect 687 -47 690 67
rect 717 -34 720 13
rect 1050 -39 1053 67
rect 1080 -26 1083 13
rect 1511 -13 1514 98
rect 1400 -16 1514 -13
rect 1541 -41 1544 80
rect 1055 -44 1544 -41
rect 1677 -49 1680 80
rect 1694 60 1697 80
rect 1711 60 1714 80
rect 692 -52 1680 -49
rect 1831 -57 1834 78
rect 1848 65 1851 80
rect 1865 62 1868 82
rect 1882 61 1885 83
rect 332 -60 1834 -57
rect 1994 -66 1997 72
rect -20 -69 1997 -66
rect -49 -84 57 -81
rect 78 -84 428 -81
rect 453 -84 765 -81
rect 790 -84 1102 -81
rect 4 -109 60 -106
rect 80 -110 121 -107
rect 361 -109 426 -106
rect 447 -110 518 -107
rect 721 -109 768 -106
rect 786 -110 846 -107
rect 1084 -109 1103 -106
rect 1122 -110 1558 -107
rect 75 -126 212 -123
rect 773 -123 775 -122
rect 217 -126 432 -123
rect 438 -126 775 -123
rect 783 -126 1118 -123
rect 853 -135 1692 -132
rect 525 -144 1846 -141
rect 1874 -146 1892 -143
rect 1874 -150 1877 -146
rect 128 -153 1877 -150
rect 1889 -150 1892 -146
rect 2010 -150 2013 71
rect 2026 54 2029 75
rect 2042 54 2045 71
rect 2058 55 2061 73
rect 1889 -153 2013 -150
rect -75 -255 -71 -167
rect 1882 -177 1885 -159
rect -4 -201 325 -198
rect -25 -255 -22 -225
rect -4 -255 -1 -201
rect 19 -210 685 -207
rect 19 -255 22 -210
rect 41 -219 1048 -216
rect 41 -255 44 -219
rect 241 -256 244 -230
rect 259 -256 262 -230
rect 278 -256 281 -237
rect 298 -256 301 -247
<< m2contact >>
rect 1067 467 1072 472
rect 1029 435 1036 440
rect 1067 424 1072 429
rect 925 382 930 387
rect 943 361 948 366
rect 1027 408 1034 413
rect 1336 420 1341 425
rect 1383 422 1388 428
rect 962 354 967 359
rect 1688 409 1693 414
rect 1701 382 1706 387
rect 703 325 708 330
rect 738 326 743 331
rect 774 325 779 330
rect 943 328 948 333
rect 1023 325 1028 330
rect 1069 324 1074 329
rect 1142 325 1147 330
rect 928 302 933 307
rect 962 303 967 308
rect 705 279 710 284
rect 736 260 741 265
rect 776 260 781 265
rect 1188 279 1193 284
rect 1069 260 1074 265
rect 1380 249 1385 254
rect 1405 249 1410 254
rect 1459 236 1464 241
rect 315 224 320 229
rect 672 224 677 229
rect 315 203 320 208
rect 672 203 677 208
rect 1032 203 1037 208
rect 1395 203 1400 208
rect 1636 168 1641 174
rect 1636 149 1641 155
rect 1789 149 1794 154
rect 1951 150 1956 156
rect 1789 131 1794 136
rect 1951 131 1956 136
rect -1 -54 4 -49
rect 356 -42 361 -37
rect 716 -39 721 -34
rect 1395 -17 1400 -12
rect 1079 -33 1085 -26
rect 1050 -44 1055 -39
rect 1559 76 1564 82
rect 687 -52 692 -47
rect 1693 55 1698 60
rect 1710 53 1715 60
rect 327 -60 332 -55
rect 1847 60 1852 65
rect 1864 55 1869 62
rect 1881 56 1886 61
rect -25 -69 -20 -64
rect -1 -110 4 -105
rect 121 -112 126 -107
rect 356 -110 361 -105
rect 518 -112 523 -107
rect 716 -110 721 -105
rect 846 -112 851 -107
rect 1079 -110 1084 -105
rect 1558 -110 1563 -105
rect 212 -127 217 -122
rect 848 -135 853 -130
rect 1692 -135 1697 -130
rect 520 -144 525 -139
rect 1846 -144 1851 -139
rect 123 -153 128 -148
rect 2025 48 2030 54
rect 2041 48 2046 54
rect 2057 49 2062 55
rect 1881 -159 1886 -154
rect -76 -167 -70 -161
rect 1881 -182 1886 -177
rect 325 -201 330 -196
rect -26 -225 -21 -220
rect 685 -210 690 -205
rect 1048 -219 1053 -214
rect 240 -230 245 -225
rect 259 -230 264 -225
rect 278 -237 283 -232
rect 298 -247 303 -242
<< metal2 >>
rect 1029 413 1034 435
rect 1068 429 1071 467
rect 1388 423 1691 426
rect -75 382 925 385
rect 1337 385 1340 420
rect 1688 414 1691 423
rect 930 382 1701 385
rect -75 -161 -71 382
rect 944 333 947 361
rect 705 284 708 325
rect 738 265 741 326
rect 776 265 779 325
rect 963 308 966 354
rect 316 208 319 224
rect 673 208 676 224
rect 213 -13 216 109
rect 569 -13 572 109
rect 930 -13 933 302
rect 1023 275 1026 325
rect 1023 272 1036 275
rect 1033 208 1036 272
rect 1071 265 1074 324
rect 1142 270 1145 325
rect 1193 279 1495 282
rect 1142 267 1399 270
rect 1395 266 1399 267
rect 1071 253 1074 260
rect 1071 250 1380 253
rect 1396 208 1399 266
rect 1410 250 1481 253
rect 1292 -13 1295 109
rect 213 -16 1395 -13
rect -25 -220 -22 -69
rect 0 -105 3 -54
rect 0 -182 3 -110
rect 123 -148 126 -112
rect 213 -122 216 -16
rect 0 -185 244 -182
rect 241 -225 244 -185
rect 327 -196 330 -60
rect 357 -105 360 -42
rect 357 -225 360 -110
rect 520 -139 523 -112
rect 687 -205 690 -52
rect 717 -105 720 -39
rect 264 -228 360 -225
rect 717 -232 720 -110
rect 848 -130 851 -112
rect 1050 -214 1053 -44
rect 1080 -105 1083 -33
rect 283 -235 720 -232
rect 1080 -242 1083 -110
rect 1461 -193 1464 236
rect 1478 -178 1481 250
rect 1492 -163 1495 279
rect 1637 155 1640 168
rect 1790 136 1793 149
rect 1952 136 1955 150
rect 1560 -105 1563 76
rect 1694 -130 1697 55
rect 1711 -163 1714 53
rect 1848 -139 1851 60
rect 1865 -163 1868 55
rect 1882 -154 1885 56
rect 2026 -163 2029 48
rect 1492 -166 2029 -163
rect 1478 -181 1881 -178
rect 2042 -178 2045 48
rect 1886 -181 2045 -178
rect 2058 -193 2061 49
rect 1461 -196 2061 -193
rect 303 -245 1083 -242
use NOT  NOT_3
timestamp 1698475750
transform 1 0 61 0 1 -100
box -7 -26 25 19
use XOR2IN  XOR2IN_0
timestamp 1698769192
transform 1 0 106 0 1 118
box -106 -118 213 101
use NOT  NOT_2
timestamp 1698475750
transform 1 0 428 0 1 -100
box -7 -26 25 19
use XOR2IN  XOR2IN_1
timestamp 1698769192
transform 1 0 463 0 1 118
box -106 -118 213 101
use NOT  NOT_1
timestamp 1698475750
transform 1 0 770 0 1 -100
box -7 -26 25 19
use XOR2IN  XOR2IN_2
timestamp 1698769192
transform 1 0 823 0 1 118
box -106 -118 213 101
use NOT  NOT_0
timestamp 1698475750
transform 1 0 1104 0 1 -100
box -7 -26 25 19
use XOR2IN  XOR2IN_3
timestamp 1698769192
transform 1 0 1186 0 1 118
box -106 -118 213 101
use AND2IN  AND2IN_0
timestamp 1698685374
transform 1 0 1528 0 1 93
box -2 -15 94 58
use AND3IN  AND3IN_0
timestamp 1698684844
transform 1 0 1678 0 1 137
box -18 -59 100 27
use AND4IN  AND4IN_1
timestamp 1698684672
transform 1 0 1832 0 1 136
box -18 -58 114 27
use AND5IN  AND5IN_0
timestamp 1698684513
transform 1 0 2008 0 1 137
box -31 -67 121 36
use NOT  NOT_7
timestamp 1698475750
transform 1 0 661 0 1 337
box -7 -26 25 19
use NOT  NOT_6
timestamp 1698475750
transform 1 0 751 0 1 337
box -7 -26 25 19
use AND4IN  AND4IN_0
timestamp 1698684672
transform 1 0 825 0 1 340
box -18 -58 114 27
use NOT  NOT_5
timestamp 1698475750
transform 1 0 1165 0 1 336
box -7 -26 25 19
use NOT  NOT_4
timestamp 1698475750
transform 1 0 1043 0 1 336
box -7 -26 25 19
use OR4IN  OR4IN_0
timestamp 1698685870
transform 1 0 1774 0 1 317
box -25 -54 100 28
use AND2IN  AND2IN_1
timestamp 1698685374
transform 1 0 912 0 1 403
box -2 -15 94 58
use NOR2IN  NOR2IN_0
timestamp 1698687859
transform 1 0 1174 0 1 466
box -25 -54 22 28
use AND2IN  AND2IN_3
timestamp 1698685374
transform 1 0 1305 0 1 436
box -2 -15 94 58
use AND2IN  AND2IN_2
timestamp 1698685374
transform 1 0 1690 0 1 398
box -2 -15 94 58
<< labels >>
rlabel metal1 1406 -15 1407 -14 1 gnd
rlabel metal1 301 354 302 355 1 vdd
rlabel metal1 1069 509 1070 510 1 voutEqual
rlabel metal1 1419 513 1420 514 1 voutLess
rlabel metal1 1626 511 1627 512 1 voutGreater
rlabel metal1 -74 -253 -73 -252 2 vinEn
rlabel metal1 -24 -253 -23 -252 1 vina0
rlabel metal1 -3 -253 -2 -252 1 vina1
rlabel metal1 20 -253 21 -252 1 vina2
rlabel metal1 42 -254 43 -253 1 vina3
rlabel metal1 242 -255 243 -254 1 vinb0
rlabel metal1 260 -255 261 -254 1 vinb1
rlabel metal1 279 -255 280 -254 1 vinb2
rlabel metal1 299 -255 300 -254 1 vinb3
<< end >>
