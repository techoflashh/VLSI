Question No 5

*temperature

.include TSMC_180nm.txt

.subckt NAND node_out nodeA nodeB vdd gnd

    Mn1 node_out nodeA node_y gnd CMOSN W = {wn1} L = {ln1}
    + AS = {5*wn1*LAMBDA} PS = {10*LAMBDA + 2*wn1} AD = {5*wn1*LAMBDA} PD = {10*LAMBDA + 2*wn1}

    Mn2 node_y nodeB gnd gnd CMOSN W = {wn2} L = {ln2}
    + AS = {5*wn2*LAMBDA} PS = {10*LAMBDA + 2*wn2} AD = {5*wn2*LAMBDA} PD = {10*LAMBDA + 2*wn2}


    Mp1 node_out nodeA vdd vdd CMOSP W = {wp1} L = {lp1}
    + AS = {5*wp1*LAMBDA} PS = {10*LAMBDA + 2*wp1} AD = {5*wp1*LAMBDA} PD = {10*LAMBDA + 2*wp1}

    Mp2 node_out nodeB vdd vdd CMOSP W = {wp2} L = {lp2}
    + AS = {5*wp2*LAMBDA} PS = {10*LAMBDA + 2*wp2} AD = {5*wp2*LAMBDA} PD = {10*LAMBDA + 2*wp2}

.ends NAND

.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd vdd gnd 'SUPPLY'

V_in_a nodeA gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)
V_in_b nodeB gnd PULSE(0 1.8 0ns 100ps 100ps 60ns 120ns)

X1 node_out nodeA nodeB vdd gnd NAND

*capacitance

.tran 1n 600n

.measure tran trise
+ TRIG v(nodeA) VAL = 'SUPPLY/2' RISE = 1
+ TARG v(node_out) VAL = 'SUPPLY/2' FALL =1

.measure tran tfall
+ TRIG v(nodeA) VAL = 'SUPPLY/2' FALL = 1
+ TARG v(node_out) VAL = 'SUPPLY/2' RISE =1

.measure tran tpd param = '(trise + tfall)/2' goal = 0 

.control
run

quit
.end
.endc